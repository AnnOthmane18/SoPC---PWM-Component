    Mac OS X            	   2  �     �                                    ATTR;���  �   �   �                  �     com.apple.TextEncoding      �   �  7com.apple.metadata:kMDLabel_6fewz4cdfdzgktx5qxtxynvksm   utf-8;134217984��Ͻ��p�\đKv�$Tyw�j#c|a�)"+|�͂�f����U��&Xq�d�����K�����c?
�<�� ����HS���jW�a"��+�c����O�c1mb~�!�1J}1��\�Գ�4x�:��%���RK����IX3|��P�a�L'j���+k�~�`LfA�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       This resource fork intentionally left blank                                                                                                                                                                                                                            ��