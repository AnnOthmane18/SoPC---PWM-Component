��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n�2uO#)�Y>�P[!W�n)6����o�hY[�ܾʰ��)�q�3����ϺeK�^)p��Hz�{%,rU���_��^�^ۜ���l��1An"3�"�����o��LV�laD=tp8F�Xx�(c���J3v����=�I��O&��2��O�j
m�ҡ��rz�z�v	R��"�R��췰Z�ʁ�����,�>�����P��$�Y��B}�R�w�Y�["3̊���e�Hʩ�D�$���s2�l*���)f�|}3���K�q s�])a�'�<7�������0ꐿ�	�O���K�"BH8>�?�ψ��ޥ���Hd�I-�m3v	G�W=U5}��JMi=���KR5��꯼p	7���{����z��) ����lʉgv���:rf�m{v��9�3�B"���Ԩ����+�p-2�9ᔚ��Ao�J�T{���i8p]E�sd:�R�����Iv��t��s���}�'��bR2m,� �Kɾ帢���N%3gv�cٮy&��"\��m�ia�J���|_�������y�����]&L�]Ш["��|�
���Pk`�e�,'8M�X��|��4��g�	;N��P�D���i6�M:Ǔ�\
Է�l7�4ݫ�ZEܧ���k+;>��j�K"���1�6�G�^Z���.a������7/��C�v�~��yz�e4:�e�v����6� ������6��B�,��`[�"	"J�E�L��SYC�|rͽ��Jqa���3��5CO�M�i�f1x��g?�O�OR��xFF�⤻�j��B�f�
�kJ���&-)O�,�g���+K�h��1S��P�=2Q���w�����y,����a��&�A"~��k��<dmg�*/��1B�>c���g!4?��d,���9.m���_�H��lz�N�6N��~�	��K�6o�`����'<���9��$V��,|�0b+���t����b�!:BNGc�-{������	.����F��N>�ʐYN#�� ��
�y�%�YQ�V�d ��V��>c�G�v��<��4ۭ�n�~��,�gxK���U'�"خ��s�(�p}��{�8/N���@�X�BԨ:i�$zy�$���2����d+;��]h��P� gz�q|b�����!`^%�ΪIw����bK�2�,�ٙ���/�?w���eՀ�m1����ʧc�g�V*.��хF�B��;�YN%�S�2��SLA��sb�V�����1#���a��3uCB��Hռmm� � ��/���8H�M��B�@�̋e�++��G6�,�KW�|��~=:8���K�$����X�T���n�3�������4�C-r6���:�B�������q� �@:�N�W��Ȫ�&�5㽮��	�qͼ��fG/��dA^�M�cg6��ʳ���2����A�l�͜s{�`Ֆ�}s�
 �^��V���
�w����À��
ûr����
Ts�(�It�q��В�;\��ٌS���|Hh@�I�K��>�r��~����(~{&lD�n���W��ϕ��Nu5IB���s�_�k�� ���i�H���!gN1JA�%�&�����M4[���[p˒�
%۳��8d����@���r�ͻaD�/q��7�{�����,��mbd[*+م�ͅN�6c��o��󟓂O�ڊy���>5�0�t�"�j�F��?փ(V�/��3T�,�vh��{?��p���Z���Հ���uI�c�����Q�P�O�4ƲÙɟ�Ѐ�ӧ�K���q)���^VD���d���?�m��Q��2����/˃���]�ڀ�z�m��Jf�F|Z
Q�p�8(0�@�kb���\u�`5r�Yj�
�o�_����"�I�w�!�{!�:�*Z�؃i�dg��a��7�9ׄw߂c�N.����x.?��*��{?R×��KS��H �K�+cK�Y�<$Y7��/H�:�|��>�V�B���.%枰���(�yN@y�	'�V�����ׁTٰ�l�xab5\x���@P��z�		L+�#p�X82��z:''ռ��v4��9�`ԹB�$=0��E�ui�]T8U��䙈�,r�T�.c������vE�3Bx��S�����56rJѓ��� 3�kT��i�R E/M�Ʀ.��x�,�����S�D���P��N�L��M�F��NS >s��s�?���A��1=��$r�af�6��R,Ȍ��"����q������Y7�}QD�e	rI���
�>�E���:��9�o}a�R�d�i�$�yǞd�K�ʨ�*����#��K��(�͔���H��Tr��+M��&��P%t�-�� ���n�r3�x%f��m�P@%�P��o�e��t*����3�9�B������<N8�f
�V�>���s
q�/��QA0��5�5L'D�s6Nq�\K3����		nm��})����;�쁩i;�G �1����E%��5v7������Ȍ�D1z�0��M͑K"���gu��;*{�g��� +�JV������7����IQ�o:�qi=N����˖�V��G^w~��ʞi�ϴ�>9��/H9 �,�P,b&�/�ߐ���8�9gǚ�-|td��#+�0�B���C�s>��]�R��B�9�i7�Jw�����K ��R�1�eL��z�>����֟bo�J:��y,A	P+��Hk#�ǧ�~Aִ
�V��7o�DUg���#>��?پ�	ǝ�c���?u�@���+�g�8�3�)�J͢��)��5��Đ-�l�B�Y�Bq�5����m+�/�r�=�-�y�s!�Ӊ� Џq��!9�I�0�V�n:ƹQd=Z�dU%Dq7���m`��k�.�A�T�����FI��n2.�m�k�	9A"D�ρ�WAU�%Z"�(��x�O!�����2n K�~,h�^W̢C�=��yr�;	O��:ـ���9�
Z����Qڹ+w�oz�Q:2�?�ʭbp����[���T0���O���7�PfFh���Jr��A��'[4�������=A�]c�M�?�rK�ߣ����oLyݽ�J2_�3��>� (&��"(�h�i>�܍�)��/���m�#�;R>԰B�	�u����y,�Ӄ^��C�����/����} r�.�NAfZgj���C�J�����^lW��E�B��*����Ng��>~��֦B#��m~I��]y�͒ml?�IX�"E�
B�N3;Lp?x%����o�ɩ!��Y����L��rKd�;$8V��yI�*��wD����=���|UNj��VD�=
�a��/\׻C��XU���L
�A�>�
d��X��m��6�TC�@Tx�\�ܩՁ'�<#9�s�Z��ύ̒O�8׷�8WD���np�ѭ�Y2�\��h?��&��t�@B+e��S�����6�S�&��+ndg���ZK����8�L�,��Z���{=E*oܿ��N[�WY5\��%2��0)�IJ�o��v�O�������|�b��ـA�ᢪx�E���1�l�f<���lQ�����¨����U�q9�x��u�)\��w��M	8H�X�����_C�:������\��/nc����5�a�P�U����^^epZ�4���Ξf�	���´B�rd���0k\Q�4�f����i�!8'G�DC��(甊. ((mL��G�s�&�)
왶��մ�v-���6��ѿ����p�6X������_����?��2�t��WY FS�x�q[��������jP����?A �
�c�y'{�3ȅ�BT�6A<!�p��E�����!�BpR`t�g7��dh�X"ρ��H����G�X�K�k�b��Y��ޜ�Zs2��7�+�KN�Gly8�,�mP�䋕����np��?��f�o������'���}��kt�u�s�~�C~�rC��?����Mi�o�M(Ԏ�9l�,��X��~+t�WL
1\voF����۪���0x�u�&;2#����!=��\1���bx`<h����m���|�?#�V��e��DVP;)�Z���+Q+��	o�0,��N䢞�>ۓ[���$^d���/~E��q�ې_oL���&AqV�A݁��d.+�^�k���lD]J	� J��X�7���{���q�C���I�=��_�*�&p�U<�6�y�c�J[�SK��1bSd�gq��<Sf��U>g�|�9ڇ쁖~�`C�At#����i(�s Ԙo�KD]����_�����m�!e�(�Ki����5� �e�6�A!,3���pE2ӑN� q�0C?����&���'��U�#4��AٗEGz�[�A�Ͼc�a=��p�?�Ӕz��G��;ᇛl�p
���цP�"���q�$��hy_��E��A�H�����t�E�k��%�����w�
�VqY���+π-���"��mzy�`Bq���^��g�T�Dn����q����4�)�0N��_�u�^���|4T���|4�&N�/�yL��Q�w�V+&�О2�<�RT4�Y��N�)4E��t3�����8a�jj��R�Wm�E%p�g�p[�U<+�ȼ���sc���t�fn�=0��=�W9�����K��6`U��U�y�s��f�[S�����������:�j\��AQevGS:�[��L�j���_ �:�9r��t�u�U�q*�t�oB��Z|��܈�~v͍鿇���LA魓w��R��tl(#�ȷ��U}hP[k4�nX�U����lLcg\���t�bG�H.�T6��~���p��񕜶�%�m,W�9��CM
�.v�U�ǈ�mS�i߭���[��lN$ʓ�M6d��֊���G��C���ۢ��[{�q��uv�J��Rݾ
�@�ox�"�*��-4�E�C�0�V���dq��Gs���ǰ-�Gsj<����6����R2]̶�<J ��s�
��i^иCK���N��t� �F��4Ǟ8Y�^O�^A` 
v"�gÙj@l�:��hʤD�g�z5�u_�5�澈U�`��n��X �6�����G�pA����OBG�Mq��:�1󥉃�����$��!�K�M��S
���M<�W}���M,�*dµ��֥�>��JotB��8�� �fu��nm�p���[���������JhQ�~�z�����Ŧo��>�Zl�����9�Ө���Y$����~ｼT��c�U\��=�k�#����{BEhv�a���|W�W�Ib��Eu�0A�5��x�eN��T\�:��,F:�E�%&��A�&.ǉ���ZLkؽS�}<��+*��ug�L�SGC� `��uR˒VϿ��";�5�f˺����Ⱦ`ޫܳr!��k+����k�f �3&��$��`ƥJ���h0���)a�!���t��n������kw�t�24 �
^�m�-8F�^.-�㗒[��Yy �掶S��x�f��
1��ES��ҟl�	H��l����ʓ�Lݘ����>��P]�Գ� �5�_.~X��U���)KWҁ=;,ZZ��چ�,2wC���<�Ӂ;,�:W�1m��U�6,nI����3�������7Ǉ���v26d0�ο��EZ��<��\���FX�=-6��pk �����絚�����.�_��TK4{�d��(��i�CS2J[�Kanj8[qɡoNew���u����� 2��I#�IR�>b�;nۄ6V�1�=9��֪�7��}a�.j'��|�B���i��Df�����S���W)�=h���E����BomBj[s(dG�ø4�C%,t \��`g��!����o��Z:@�f��������𛮑:�#�p�}��: p�		��yI��m��\��6�P�m�,{^ƻ8���5	P.�1ZV�h$&�u��z�Z��%8��KM���~�|��5/�z�B�m�-�z��"E-�����
S�7�e������)<C'3<Z�|0�% F�Ֆ��n�ؐ������;{��w�$^�̽������eݙ8�|�ɒ*��rɴ���1Q��A�5"	`�t���\bZ�W/U��ׂ���M����wU�����8'.����2#y�Ӂp�V	��sS�uU��I3�F8?�n�<yy�K��74�	�|�=ݷ)iA�S�ec�I{v�kB�|��G����0 M�X�9��EDG�Wd��\~9��Jj4���!>��)5�����pU';=�Ղ�:�|�	mm�A�Dqu���l�����'��=�?�2�ʬD=�l?s�>�.� %A��섭���u����@�56Z(X�7ȳ������)f'�A?˒ķ��?�q��`���M�h� ���Y"�Q̒�����M�O��4�4���j/,���r�\1� ���qw7.�����x�rl�O*/�9Z�Dind!��_)�X2���� �x�"��O�6/ץ�m�/�WQ�~��I-�B��Hܷ�h����[N�G��`+i�KB73�+'�Aчº�fR3��@���IJM��Q�	�����E`q��{;~)�Z�߶{fW�7طB����dp�g�j�<u4 ��;ۿG��Y�����GbQ�FiF�<�8X��XD�f��j���-��1(�������J(TD�N#ǩ���<)Uή��ц`���at�k�]���bЋE�c�U ���hmc��%ݜ�ɢ�)�f�%�Z��W��H�r�|ic>ڢ�:�/M��e�{ZӘ-W��m��8��[�F��\��U����N�룖���&��g.'(���$� ���0��] �HD���%�}�9/.��!�hjɶ�tK0Y}��1�l��Z�kߏ�v��4&0���tʯ4��JyT┤ݬ�v���bfW`Lz^L�:�1�^q�rncSn��gO�u�׆�u0�x?�ab���d�q��S�xPܙ9��Z4~VrT�ۤ�����n�Q�ثx�c7�kJ��Y���H�C�o"]��)���i��{��:���"�8��
�\o�����L kL�_Ň6$�y���ư+̹�����k1d�\�+p��,�d�E�Qp;����F)������M�z_�P�`��l���[�u=rM��h�&���:�nt����H&��=�8+L��ႜ
�Ȼ���36���G�<��>��*:�h�yx;����C��\g���c�h���w���?� 98WAK0�\�[�av,�~��WT�Yn�!���1K����%[&�&9���/�bʪn�*#��+��5��D�4����K�����!��;=��������9�	�N��<űp,H��dk9�m��]���5�ł'�_�uaw?�Yp���N��f+�c��{��$�n��}�%�Bo	�W�jѕ_l63���v^� ��j������;x�K�̠���ބ.�(zjˎ~�l*�wV_� s��Vs�Ss��C�T�.%:�9����Հ{ʌ�0Rf��R)�|�3��~+ {2��LxW��=��S4<a����p�j�޼�j*�c�]���ߊ����wk�9����2f��.Фw8@�M�hr-%�>ȭ����e���L;�- ��F���R����ܡ���T3:U�f�z�8$A"�k5�k��`�&L��҃�9��UL)�S���,�%)"|ΗꐫXs0�8$e����R�I�(S� Pp�-Ў��Z��]��b*i^�&�$o���")�5����#D���J��)^���^F�ߍ��wR�f�F��O,
�U�n ������LZ�y]/�Ϡ��K�f���n��"���dP�ދ|s���K8,��n�&��4�.7�~̢�%���{�EfU��Q39�l9�-��ؚ�d�h2�]�.��@�S��!?�O���c]�X�8�?�;y<�S�ng����.�>"��`E��Ʀ�EZ��Ue�b6���ͣ�A&��`�`%���¥70��wB&���T
M��� qU��z�W�*$b�=I>P�q5��H�Hǈb�����p^���߿��;Z#�i8���@��T�n�Kb����7{i�F�+�'J�*�3��^������dtI��a�%H��l��:m��%?�P]�"�$�(�g��:����6��<�ɜ+��d2	1d{Ė?���d��aY+�/7x(n$�[��ŗ�5c)��!����������z~�=���_�A!D=8Ӝt����dd�deRԃJ��E ^~��gH^?��GX����Y}��K+|Ր<�n7�z��?�	!���Į���g��|�k�:1��zױ7�=H���F��~k[��{Է^B��������b��TlL�b��֑���bW���I؍$��)��2�����Z�i�5~񩥯3���_�?w�j�})��C֙K��'�V�]
�on1�y��x�#��{'ڐ��5�_��� �9OT�֐��;�M�讗�RG��#ߒ ٳ�*��ˬnt�G�)�S����l����-��Bf�n�E+�M>��H�j����CJߟڲ2�+T��̌ ���ml��	l�O��3��A�6(3?����i(~^,����VN��L��?|C�3�� �|4�>�����0]d"8{���\���Y�J��F��%z��_S����U�9	��maK��^޿R��Dc�m����/�ZWat��k��}��i"�P;	o�e+�)-T@�Nyӷ��`�O/~񻳜H�lݻ�ʃ2`�i'�^�U;^^]��ҡRX.���^]�]�v:���|5���s�'��"�D����Cc���g��-gob����c���D�RLb(���$sӡ"|L���g���r��}�	'��$�C���D�a^��g�,���>�N��"�������[_3��UI 2�"� �=�մF����R��>�f�{Y?�'-���qgifks=m� �-ڵ2Vå�K�n���� �3���yP��B�k4y����b�}�י�N͟U"N�!�5�П0'�%�A�;���Z�5�m���&�@[��<���X�y�T�iGw:3YE>�R�R�D���ˮ̣&^�U�D �CF?p(�3��2�?K}�)�:�
��m�a�b$V'�����ۦ�:ۿv�/ɏ�Q�9�+�͘޹�}tM߹_�X�U^��Q:1^f��]&��u���k���gy>7���T�g��sUh|fg�e���{P��,�5���e߀qQ[�1n_��6g�A�m��%��n�P�<oxOD"�w�2<ۏ�~�~g��+�;�@��;�Ǹ_���C�xo����ؽ��Yt��`lGZd����"�ʴ����y�6�Nɻ�j��W����Wj�Z�}��g2P%�xU�+I<�j=�� �1�)��
wʲ��`<N;]�no�?ɓO��Yy d gi���i��*�-��-�:(72|�����u$&�Q/2���_ك��j.�5�!�o}�#�c�t`;,�E}���_(����]�ƴ�AtKo���[�@Syr��b�n3�F?afj����� ��Ƞ["9�s}�s�}�0~����,���y<����_L�-�Yb�q7�g�(�+≻Dil泓�J�������n�U�{yE+�Esi��\���D4�_ʋ>���^�+���w�C�o�f�4��
a����[��8e�*�^f�ǲ�0���l�W�=���ۀl�9+�F�E`=�� vJ]�X�	���y?�?_������d�
��Ӽ
��D���fW'C�?�rP6�^N#Հy^7�VK��,�1Ku^�T3[���}�L�k�4H�|̙A ��s <s�2So�]}�%}�2�N���[�E�$H�$��b1�+k~d�ہ\��m|jd��'3���0�s�qH��+~"�W�R�Ћ,[�WY�枳 �	�4����H%#n(<G-��������}SP��R��m���5.l:d����maa�%Fb�Kd����'O�_��g8���;KɟU,�0��S�		MO%��D�A�m~6PpS�B��ΖRr��^x,Pn9f��LgY�]��zܭ�q��_����	�<N��#�.�eS�J����I�*3�g��>���þ��o�"n�E/pf7�΅i�����^ۺ���;��b�wqlw[bPJ��<%Z�P�X��L��,�J��&
��* %/e�zv!�p�O[��@��J�9Q�a���j|�d~������(*�0����V�^A�HUS�aҕ��[	���{Y�@����J-. �!�0��_�hs;�Q��A���
$��\�8v`�
\�Rڠ%lN�j
t�,EN�k�K�q��=�)pA�[�N�1�ڊ0��K*zv^�/?���;K���KԈ�.z��L�X�L�ߜݱ�BY0���|&��,̺dX����5%zr#J�S��?�c�|%B�M�5�c�Yތ��%Am�RNk�y��Hl|�%�������q�� Q�֭�7в���Qq�t�l�1�C7�g�����a�s�A���ރ�d%e��+AL�rH��CL�j��/�6y`a93я��{9�'T?wQ���v� �^�����X��Z9��3�I�dI����|�p��#�|.�!|.1����,�(%�����>e>^�/@W<Ay��y3��]{�v��t�,y0�UcՄ�H@L�w�;Q�&����0u��}gv&5h{�Q؇���'��y?�W����	b�_r��s�h���_�{�~�q ��1N)�j�mD��2�𔮞w�h�Xk��;�Ŧ����V�.e�1e�_�~��i��_������[� ��{�t%��my2D{��Ѹ��I|"vj����AZ	S��:��|�W=T���'
�w����J} J�!Op�s5l�?��b��������I\q[|��3�ɶ/v�Ov8h�GX6&/�Q�P�ӡUU&j��`�E�=����#��aC��Yo#�����A�>��{���������=�9���S$���f�0��q���$�ƺ�X�~=���eOB�x����Z��4$;����F��l&O�������LӚ��mZw�-�(,L�餸�(� ��L�`Z9f�))�	�:b�}48ZM.���i�L�a���&���`��7)�b�q� V��tY �;X��`���?,d�<�6P�W0(����r~�^`{�+V�w�1������ܬ5ɦ�i�#���d�
EzZv��?���y���$�\�6V���k9U��a-5i��GMW)/�A�;���I�c�*���ً�^���>��T�[wt�%��n����>�����~��p`P�����9�%m����WE�=.u�C(nYM3gXa��2o��]W:y�NO�����t%W�O3�ȗ������:s�8�A�?Sa��ӱcB|>��D����7	��^��*��X|/�b��z�᱾�.�5����AvY7�����q�&��/~g�M��5��~ٱ����hg�$�3�D��ST�e�#�v�����>�=j�&p^.�Ŀ�AC٧��̶h�K~��&���!l�@����1������G{z+���J�20�"g�E�'(��x�D��	td$�-�	��"�
$l@�ZПva^$+L<������:j�ÔG��� d!��&���oԷ��68"iz�����dh���p�2��يh�Fd��شm�L;���f���v�H}jD���g٤�ﶰ�0d�j��d��L����]����N����ū��!Rp�X}'ܞ�Aڣ��|!E ܸĵ��P|��
�Gk�&`n�����X�����Cp':�^���)�F�O�(_}�A4���Iꄃ)��]x�?ό]��"g�#���*ӋM���U�������`a�wg�J0bAn�VJ�qYu\9Q~9�G�ͤ�� x8}!sI������P�{����"����_��2,YjQl e�B�4�N�W�B&)Q3io�r��R�p��;�i�
�&we���:�1�z�8g(e�)hS�~o
�]}K�s�`���v�aXrh��Z�E���WL�7�W�*����~�ru�d�>���9C`�
��Q�N]��G��Fp��Xt���m:2�ȿ���˳��2� ��t�bV���"A�T�i�m
�kp��9(����+���F�@���כ�ř��o�"��膅�6��*�Vf� Hƍ����<1�)��6�VY���W�ui�e�B�$�����$�[`��38P4u*�Y�X���۬��`j�,�䏦�8�9��˩���U;7�R���z��$�c�m�bZ9�$=�[����_K�I���B���w⸴��Z(�:�Q ��@A�%�L���Q���Ɨur�)8�5j���5:�>:��;ؤ�[�L��B����2���T�����nN�=�M%$NgO��k��s#>K��&�10�Y'�� ��8��9:��#���׹����'��e�n��i � ��m���
aN�7s��u��]ON�����/��k���K���F!o�rc�8T�<#W��I�hԛI�T#�пcRa55!{e�Mr�gz���\v�0��
�����5��p���� S�<@�F�ynI��Ɣ�q��t\�R�$��u�P�0�3c+���ס�`�xo!��?W%r8�W�^D�c�|��a��jK��-'�#ݻi�6o�5~+���1*�Vc�H��ZI��d씸*�maQM�C[P�V�V��Ԣ�$���_Y��rͫ��N�6��O�=۰
,��u;�aI�T�vk�(e�&p����ʳ��G�
c�5�k;+l�	G�P���Z"�/�z׾�+:/�Axw -2�kH��/}�V����D��-���Q��d��D1.����* ���ĚC��38�>� 2%s%��rbF�T�CBu��M����]�(�rF��${p/r'˲�O ����-����)�h|u=s�&O6�'ۦ���?*�κ�2��1�׊�
��'(K�dZK8!�D,������(˥��%.��ůpY���ˑ��V�6s�<����=��r�BW5���N� ����Jx���6�c�"�� }d��.�iQ��sq�Q����N�VIL`]+��0)�'�mQ�#V���B��5~��~r����*���?YY2Y~r�'D���`�oP�v�4��$�-�:�E������VI;0�N��S��w4�6�_x17�,TO��G�o1{̩������5e���zZ�ȷ�R�����v�4;��W��s�54����|�N��c�@�#r �a���@Gg�d;�%��nC�Yڋ�4Qwlu5cG]�k�(��,T��_���b�p?0����<�ƍ�g����D��N����T�hĆ�P꭛�����؇;Uw�D,�ZY��ŞG���Ix��Y���%Hov���?����Ep�@BYk,�/k��ܳ6� �_�u�P�|p8�o���t���f{���o,�}X/��)��{\b�kN�"�U��	���|��"r�y��
�����u�0��a��T�R���C�-��W���g��sq�]�H��w� *���I�4Q��.���)��\*k!�&1I�D��u����KǤB��L���ؾ�
\��S�&�~��N���쳠�MN[�R2��+��ltN�拺����J����
����F-m9��B�mo�����6�NH�WS@6۾��1�Ρ��$�� 
ިܴE�t�	@��>�Ő< ۇ�y�Zs�� /�ݳ)e jn���:yi�Y�1��_�ސ3�Ʊ�F0������[�c�z�<{O�:����SG�[7��2C���M�̻��� ֜ #B���ou�*�G���V����>����S6�-[��@-��h�%s��de�t��eϳA�_��-#�+�~�e�3���+�9?��\�y-o�\������cۧF�+Epq��R<�Rjf�L�F9+~��C���Á�={��y�?���a�^��pbj~�a:K�3�ԭ-��/����f���F�x2��KnCͬo1�5 T��*��c���i�GD/��N�:��g�
L���������xN���!�B)��}r0ؙ_J跍�A#}C9c�m5��#X!GQ������xh����|�6�#<tYn%t{7��7,cя���(���w&Ⱥ����y���zfBs ���P�)~�l<T �⨙��9�V(���b��H�ȫ���RG�� ��\�Y~ט����߼]��tE�|A(��0ƛ('3f��ɥ+h/L/�6X�9�>�IF�{5�0�U-e7t�,A�n	Bf�9<b8"����N���)��A���5jؽE����np/������@i`T�F��|Fu]�+h�N�>�� ��;K�k��y�Ʉ˪�52+�{�;B�{�*��4�`����33�.��l��&�@���"�ޕ���/㮨c]Paq��]^ �Gaa+�CK{�NY��h�Y�IL
�����|:��B��ސ�����籥��Y`V�Ҟ.��~j�1���J���������h�Y�$�^�L-��ʯu�h1��{R'�l������i����)y���d�S�:��F�(�^0�p�ad�mG���SyLn���`���g��h0�>賠����+%�H��� �����=k9W^�x[eD�+QR��2��Ѕ߮��L�(M4g��	�Ll�?��k��?�o��@_���v� {u6h8OF 9S�7�}b���ϺPN��t��H�B�3L���S!���ֻْ3M�t��J��O`|��Ƒ��Y�K��	�;<�|��8kO���0��/�'��S�������}���㒧��躅h�)W+	�h�\���:�bO{�rXX%���G[2,hA�����B�~��2�����esF�|�����ٕ1�U����^�	�pbW�
� R�n7��n��Q�0=�nb�G�."*�TM#!�y���X�n�a��w���3xSSwӛC32�ͦ6���)���J��7N*�~���J��yrw�)�뉈�Q��
��;�OEօ/��qlX#�E }�`��S(�7ٜ�&_�'o>�2'��n���On�y���/��ݎ��D��7O �ZcX0�t�2NF%y�{���`M�˟\%|=�HG���Tw���D����;�F�o#�����#i��U�Z�++���*}&�4���/�l�4����&�Q�,��gM������ ���5b�d7�#�P�c�7�hؘ'�k�����v�����V�RB���LC�+�?s+������� Jc.yb(��5�3U�'�4���m����ks*#W�,�h���zu�c�����hs�kGV+uݎ?�#!Z+
f��s/h�D&4n��t��p1�y^�H�K!�E\��ft�E���P~�i�A�qV�����������É���m	�-?*{_=�����v^O���Ɠ�`�Du�j�2�Qt������&�I�c�7�$!,�OҢ�84����σ�ݱ�Ů�&�y�~lP���P�q��a'n��|��œ���Fߵ9Q����1U�rޜ��S�p�}�kȣ�i
��%�	�2�Ab*ݯ�1��Mn��Q�Ц��R��T\U�.Z �X�T��!�K繚�f��n�hJ��2_a�ȼ+�	�E\П	��܎��|f��Z�E(8wa_�E3�muA�韠"��h�YP��H��lL�&!71��J�^�G�7nWУ�1NI�g"�'�+�6�������ǼFe�0�l�iK��j�n� j�M2�38�S���A�YϸU��<��`\=�p�
��B�c����[n�+��-���9��R:��F��m�գ��+ã	)�h
�GEH�l{
u!E�k�yG�`w�A1��EgO�$�T�RӮ@�{I֦;�3l���Ӽ�X��&dG��a$�d��x�a_	�(ΰ�w�Ll8�=�'�M�����h�o�ұ
W+�@%����*�O�n���ٵ���6~�۰
u>�T���?kB���V���x� �$Ns����2X�����\���{���I��ۊЅr��4 ��k�vC(�e�)3��	�������B�����A���'[��%� ��޼C�qՕ��?}��F� ��j�N��x!Q�?�58�}ޟa�L� ��z�����#��ί�;Ї9�S'm����r�ν=��Aih(m��������w��B��!p�c��PR�����:���J�H�KJRtۣ�rU<k��!�a��Z�^0��i{�{S����{���p$�^8Ϧ=�����7��sis�)lAx�E%]�1S<ܕ��!
��J��C�E�����OG}�1w���ֻ�\�d䎫���Ovhn���1���	U=���b�ׅNڶA!/~A����Kb���qWX$��p���F��d�.aJ[�C
��]�d�ލ�/�U]�meAN;l��* ����x2E�4ȡ��w�~��(:�����o%��|�fߖo�Z��ׄY`$	�O�j7e*�+�-�S1@j�i�Q@�\�:�������Ӝ���)y0�Y����-Q�Մ��H�>Է��y�ʐ3�oE'J ����)M�m�->�)��{nAym��7�������A��)'�E� ;��N�3Pߊ?��~�p�$�F����OU�����X�C��X>%2�2�n�ī���X��75�2�,P�`e ��R��J8c�M�:GRUQcs@U�,��p��`�������>IF�O;�rю��u������"��x��lb���8@�]M~��� ��A�&.a�jV�s��a"��k��l���O������#��(��Ř5�h_�[�A������h�1�7Bp��݌�� ����ȱ�}[0{�X]�1��
�
�g4����}������.cwNdpЌ�1/ٕ�Z��SL���aC�/��Ĝ�9.�]9L�]x��j�?}�OC��Y'����|��?�y8q%.y%�r�nXZ���)�2:Mm]����]۽z���l����J�V�[K� �B�����``���juߧ�� ���s偊`���n�Pf4`SO��la���^j��(v��֙HYM:��4h�T_���ÇR��%5����
��6�F�eG��}��^1�̨24���ȍ���y���ĕ3�izC����J�$�Sp�5>˧�-t0��T�/�5����$�KKѳ��8��_B�2�,��㤟��Ru3�i�E�[:�"������<�^u�뒈E
��"H6�,4�}���0�g:�ns�p�q£�v�2W�u�u��<�O�&�>%�����Ӏ&+�7J�2�O{讗�#Eo�o�,\D��4���� �	���eH0�!<>|����Xѯ����֮�!m��ӦaG�?.x� :OO�K���u�q~)2�m������I�a��~�X������E�9)�Ǔf��R!0��2������ `��W!���Ǩ���		x�/Z��yO7���[*1�:�����&�0���E#���և�u�٭ᯇ�h8��{���`k^�0�~Q��B*�C����(�f� ١�h�	RG�L04s���8}�m�8��"	�JB� K��'s�k��ՄYn�U�~I#�z��`���h�'�GFJ�͜ۃ��UG53|����܁�;0���`���=�%��⒣gh��� �t�KH�sW}�ZS�<�cy�XVH�@0�n&md�i٬4u�#@�<�$5��6r4�� 3�srH����c�H �h���ў������|�۞j�~��3%g�y��.Q����>�oF�$1�1�(�2�>Pv/'�lRk��ԝZ��H�jJ�9}m�/�!���vJ��!6�4`��/�w_���7m�*_7�8�(�]<���*���]95Aj�� c�� [���:�m��~�n����S�%�����Ne�y�E�R�*��r�\���H�F窗�O��r���aD^,�����~#,p�*t�C��Q5�L1yS,��7t���xݷ�7��H)�62����r�3
�c)q{`�笰�Q��]�L�L����RPj���0j;�MC�_\qZ��@?*���"#�G�����]�kx�4i�G�F�12q��N� y���(�s��{9q��Ưqyb\听�aw��b������ɒ�@|�ț�I�p_M�F��Kqfz^a8d��F�-�y?����;�u���U[�?�l�IznV���(n���'�����M��vn���yAΨ�g\�}N�{'�¿a��������ł��B֙7���{�x����Z��8�r]��K�C���7N�� ��nX[�G��/�&�Ȅ^
}S��"Pr�Z�d�%�]����	�è�T]
�P�<���h'*'݆ʌ�_�g�{|��k�����7ajq�;���9�@U��%��R���a�<dR;��~U�)"�<|J���;Γ� �'��fE��n���.v�u��oGnln��R�+|A yn�"�>@�;�@Pm���o�r�%Ӯ��L�+՛L/�
��EU��]uӌ�X�L���B��aP��_O0W#��U:�Ԯ���Wϻ#3��e��H��v��_���Ud�긏�^�8�u����� ����!�E���Bh1��V�3`A�>�W�6�yp{��3ت�����F�C'�=�`e�@F�}����t͓rj&��	���z�d,�	��;�?���w��Cn(Cev�D�\��c	X��:��6���ߨ�ZPov+۞l�uCk^�NhR�����ǟ��ז:����� ��W!ShH��Y��:B2��@��Gꯁ���W	R�I�����O+t��I�يӛ�G��9�iɽϙ\�z�;^�c�Ic�p��`�{?.�8.��+J`���L���L(�����	$�n��y1&�Wm�AX{���S�b���v, ������y?�����d}$�"G�A��!����A�7jf/>tL��ܭw�q	�SPq�T�3��ܱ�^>����J�`'�a���"u���FF�'m�[j|`�aΡ��g��|��e^F��x�%>ZTHj�_�\�*��Ӭw7c�J���?�&:iڜ�E#\a�xc�?��1��"걘Ԉ��W��T.m
Wcf�l���T�?KH��1�4ڷ#�م�P�~WX"V���d��W��F4�$/E�_�ykǏbv��G�3�aq�N�~'�B��)�ʓ��a--��0=x�L�z��#��=7x,�����E0�ܚ�ӢDp��=�YQ��C{�����/��M#4{�|{��P^o]��2މ�Ci�Z&�WU�Uc6[�1�/F&0 ���=��=	w/������#�"?{�*��SE<�۟�Y���G��ϲ���ڡ(\�t	!u��YS���S��C�R7�#���vKN�26�[�9`��1c�8ϲ�Kz9(�~6C�Y�Z��w� ��� ��=��Wے3!�8�Ed��������*q�^��h��ևi��1���1�J�ڎ+CJs�Nî)ũ�9%�X-=3u�W����>郏����p�*2���t�o�%�P������e�V]S�������6�&�%L&�@�Bpg���,*d s�n�掲*L�mD��z9�Œ�~�^=n��j����[��g��i�8Ud5w+r?���"�{n@u�B�ZQ�Ǳ��Ρ)G��>5�d;Gя[��A�Aj�6ڣT�{�|αe���uG	k�k'��JOTdY�z��ؙMVP��z_N�����$AfU(~��t��!u�J_$o��#���P|+=ӮW6��e�A���){ą�c$l@�P	��s����:N�0iN����z���ω��R�ѫ�$� ^ ��qȢ��z5�MYL��'��[���ka0Mt����,b����S�%#huz�.�o�6 Sg_��5�& �F�'3h���t.����(Ll,��&N�.��XCE�T^�T��d��ө*�sI2��h��g�Y{'��@R�NYz�K�TX%c��`��l�*B�������b��4�A���-�6�h����-,ߗ���V��b��1:5�=AN���eH,Õ��1�5�J	*dܩ��B̏ ��^:W�� \�q��")l}v>�
S���2��rNF4l�z�pR�[ی���W�,%3o��D>��8V�X����V)ws�`���O���箟$�'*�����突[�ﴊ3�`��B��1,�Q��Z�[�c�'-ݧlNo	]�L�I�*�x�R��"$�!~�#{R�z�� �c��u�5���c�̅��2�_�A`�/���R8r&+�;�Ha��Eit�L�&�KȐ�^2@P1L����R"���h��>��d�WH� �*J�K�k/���.c�!���.�d��6�K�̥Y��-n���|����&�Z�%EQv��*�Fh�i��s�4�1 >s������P����U�V�u�x[g}���� [l,����b��]h��:̩U�t��|��K�k�����Bہ>Q��f1K+ ����;tV��Bo/i�Q��P�Mjx��?�t	u���?�l=�r�ߠB�{�楩�S�c;��%&�.>��hv�u��y�&)7�퀟p�
���%��-|�ߞZQ5��=K�b����ͽ$9���+�r�NU���I�"[y�U�����M�j�/����VS:�op����Xu �%R"	�Z�;�Y���=���a�`��K�J� �gK�����C(J?�����7��*,�o7����4b.�P�۷=Ћ"��ަ	r��f���~Y�ժR&��h�����)G����_h#�����r6�,K�#y�x!�������|)���}{�����\���7>��\7ߢ�'P\���dF��{�8��(�T��MR�N0F	�)6)��W�:��(:����8���䝉�WQ2�:4�ȵe��:�g�U�����"M#�1U�PW�/��A�Q��˪:����I��<�(�2NL�|��#�� :�ؙ��.
�2��gK��nŉb���P|�Γv��Tw���Иbv�?QC�}v̎���I�9mӄ�$������l�9��d��]��ߌ�|�Q��2�L˻u���V'-�s|N�i���q�I~
J�GC�A��^�L�{4^ɶ�VF��O��1�M��LF�E��(8����,A/h�8��^27��2�SH���%L�[�i���T�p��K)T�A0�P4�+9P��$P
���f~��v?��aAy>^?�w�?��)-(;q�����s�4|(9jF*�q�²��C'��nG�����"ߜ�,v3wq�!o$\��d����Mlƪd+�&D��⢐`~�V�]�� _ᖋZ�o+�a��֯K�wa�c/|Hxwv�3D��a�MW��L��8Z�XiX0ܦ���&ɖ�@�u�ƾ������^/�α&�� �q��&���r1�mt�uw�;�%AUm��B�����#�.&+��'��h��h���m������8*�`�9|L|ɘS,d��k8����<�HL�3�vr]�u�Cg�1��S5���\B��f&�	�U]A�6C(�.WeC�J��NuM���	㼎��s�HO<dg���nԾ/X��O��0V���ҡ�����-�@��Ĺ�=�7�i@���g��<0�Gvχ ���@������\�&{�a�mQB��#>��ATQf�^���,�������:�pؙ� ��B=���>!�a>��Cmq��PE���n���]��\�m�K���7eFOQJ����9��g(>�=�3ǸA*�j�H:E��Mq��
�.Q��$,�M��e�˟��M�{��)z��|�q�E�W�h�*�T�)�K�$������)e��,:�(��|��q`ĵ��<Bo{�W��G5!��4H,�qbk�ۣ;�Cޱ�����Bo��M��R۵3�'�&�
�W�?����|c�?+c��8幬-EO�Ps���,I`���� %i��=�j�RV��䘲���Pm;X����V����?�A�NH&L�λN��	�#	� u~)��ËB����wA���?r���q	�C�D�S���pN]@$X���5���;��{�����'�59<��-/��E���=�Ġ�Ma�,�pҮ?�il��Hd/~�D*a�,3���?lh������
��C�M0�aKޛ�7�1q#�)���k	�,=5�`�Pi�oX��e�����9�5���8# Y #���i�'�V�zM�%j��;���\&��m�`g���_ë������DJB�~~��)~����0�A����"y�4�#�TKH�o���,�VT����l�h8_�Ow�!"�J\p�	���`����"���tm�r�&�f[�w��u��wuPV���1�ClP|�\�L�S�V�RbN���S��][y�~���p1��L�~���6�(�~a�tc�Ý� DZ�Ҁ^<fWf�a)'���J�]�J_�9���O�F�!� ׉�dǰ�w�f����kZc~�+k
��#x��/K��h�J	�l��mo�W�L��T��#�0'��49��ºFuXi�B��<�>�yH���c��}4�A��/%��L�g�"�:hr�Rػߋ��fD <Cʍ��(C���Ӫ1��R�uԌ-ِ��^��Vxv�j��0'���s6�)�/�N͸F�?ttR�uAiK!�N�`5�i��[��N���܂]9w���N��JM꿱Y���|@L�=k��f�:窺�����iof�6�½�N�8uO���S�����&m'�()O!�-�=1MH���Y�g��?�z��l�{��4��]�<S;�U�����+�3��p	��L�[�5�y�[~!��٠���z�1�EN#��昁C��D��"}j�K�lj�t��%���G���C(M�g�A��y�zߧ�U������b�4�{���T�O��05��X�^��٦�F� x9\�I�v���#��jk<���V�'����K.Z�r跪zp��C�vtn8�,N�]%����W0t���iX�,q���:93!�P�^�DR�#&�˿��	��$����AT5�Q��;x�,@����)v=>c��U�'��wY���
�,��)Pwe�/�*����3\O;��&�D��>b�5V�Ʒ��x$MÙ�#+j >Y�a�Ϝ�A��A4ya��� �/J+ow��9^��C�kv~��*wGlc��F�$Ӳ�V!�ޝc?tKd�W���BC�C_���}�{�)�9$}�)S3�ă�d��w�q��A��6�0h����&쨸/�7s��f��aH�c|4����s
��0u��6��k���섳�����P�Ω?�&�����@9��H�9���e6ڦ'%5��:��[�Z�vCj��וbw0�f<�_�X�xW�:���  y��R�]"%��3`b9q��j�a�d/h��+>lR���0MW�YKâ=[��/==�����e�=��W��c��S
��;%�Y���I�a��8|�����|H=h�?z����ǲG��v��*햚(|L0V��b��+[2�șnA�M�'�#n���h�a�¿���?��w��s�ٰ����0��݇U���I)�3��Ap���Ƶ(�>��^#@s۱�m�MN���WE\�N�Hҍ�ڄ=�Ѻ��@�ϝu,ְ�mH�j�%O�]���Q��c�i�U��qj/��b���6zr3D�^�F�΁r<�6S�Jn��d�����O�{O{b��Q;$���Kj�g�h���h�.�Tm��ޗ�~fKT^�����R����s=NgP��ܷ1|M�}��~�q�p�wv��46�Gi$��u�-Sw��H�c��Ӷ�PO}
wO=*�<Ex��O/Y��d���+�Fɦ.-|��� ��P�C1��E��C(���Q��7%���	��m������H>w��t���u(w��ɳ��+�Ue���-�"�\�|������A �.i�<�@+Yr<".2n&qEI冫�^ڞͣ����V���ʑv'J� 5�v3D��|��{�.8��P� 2m;�N��i�4GZ5��.j�NP�8_3�Q��2U�p�$=��DE�Qc$�,g� 4�k�K���3|�=�w
w1@d�$�������<�o�WW_�������	xa�Y�V�ҋ �\���ɖ@q��(�S6���r��DW��c��_�m�� Q���=�p4#�\F��R	��^7E
�=v�OVq����d}��(�ȿ�����U�$8�����Z�֖�H�:"�8@�H�>q:�+�#�aY���e�P�����Lx�E�-
��M�㞠L���t�������	2w|���H��o� [�G����ǻ"/��Ȩ��m��v��۞I�V��z�tF��� ����t��G5��5\���FM;؟�4U�)�g�}������l��	zK�W�4\�����b˥rM��k B,uD�m_[w��<2���l���Ǿ/�ɦeM%7�1/	��5d���>���5�4AS��-��/�V����H<����ڔ�s{���4�z0~	֢���'Ýĸ�#6�w�F�'5ZΝ�!l�S��Cv9�6����a�/x�J!�[�ս.: t��\Ҳ��"���\��<�:���L~xM5�%R�jY
��"QV!�����ߪy���Ѩ�6	�$��T��D껟L�p��I��L0��'�(���)�LvG�4��=!�F	�,�;%�&���_�ǮS��2�X��?{1��ʘ��hR�KTi!�O��P�.�||�1ξ��܇T$�a�zC)�(�����m�y��.~�6s].�C�VL�Bku��9#uoj?x�شx6ja:l��WL�#���Ǵd9uk&4�;K�E�aѵ���U/��ݵ�q�\� �|L9L��^���G�"Re�{����h"O�Ǣ�������Q��a�K?�*_'�J0cN�K��H��'Q�V2@.%�B>���r)p��S�f��4���~ӌ0���R�U��b�H&6�c|C�Ə���7i�Yl�i�ZÕ��O�`mZ�7NTA��ۍ���\���p������
Ҟ�1Jq!��l��M���u["�ߞ*6]���,�E[����F�
e��<!�&���p+�j�������l1K�#1J�)��+�8_��C/��@����{�S��������Kgh���*��@|��%y	����9X���,�	��\�:���.��D�6/'�����,�Ge���$}m�9��\�o�N�v�I�K&�g!!�2XW�ϥ��s��y42`2�t���*��=���M.9,N�D=Uh?�ق�R���:�K���|"-��rƨ=ʴ�ZZ��M���W6���2K���l}=B��s���D����{��5y�U���٠+�&�ԋ��f4���jԮ�Rߦ���*a(O���M����j=Z�e%�h��Z�3�g�ʲ��{���-]��4P=cpR���d/���1R��,�J�2��V�o�$Y���X����鲉�8����f��c���[����%���#�0��,]+8�*�������ø��0L@1�
�L�ķ@��Ȫ�"�� �KC�<�����|T
�gaw����6��k�\���A	Y�N�sɐ�"�o �������P\��g������H��E7gB�>�X��*��@}���U'n�bsI�JAWe!*��>�\�
ZG��;_�T��O!Ŕ���;W&���Rh�1���2r]���j�i��q�4,�i4?��\�fg�ơ`�9�(��a2�[Z�}��$+��f�Bp���,Cww	�4*�{e|4�Q�,�SÉ'�?��}@a�s5A����+�\���j�G�D�I�0��9H)IWX4�Gz�E��w^����m�`da[h�B�^ {�p��AY1�f�3��pgs �N��q����|��G�q! ����lϏ�i���'m��;2pob�es��C{� �����W�8���f�����ו;M����ð�%ЊC�}��ԅ_Q����jܭ��S����&gU�D-짉��k��������2��i?�-��«<�*]}j0����O�>�-z��8L���Q�`A��a��*^�h��N��!W-�s?nZ��ū5�8��i��3[�"����<_�x�h�p�6?6�G�4����ŷ��ⷙD_p��PZۮ�M�'K1����'�t|y}%�Fg����G����@��q����(<�b�S:����$��͝��O!�j�x�#9_�m� ����R8��%�2
���x)���I�ʓ��ee�����7R�ph�g�`���E�PLs{α���וk��T@� Zb���vF��*#�ui�bS|��O\6��^�1���1N�z�����D��3���@�Ǧ$+/�������^���8��g�]����D��o���d�!��g�7��d+�� �.m�8�/��Ӄ$#f hU��6m�w���9�ĉ��f���9�U}��e��w�aK9d1.ny���0���4?�Dpv�1�l�*n"$m��Td!p��/�F2[;��?�i�M�p�O ���^D�'R,�)�pt�vЀ?g���P(�Wb��f2Iv؃@���ZU��
���u�����ŨXi��c�-�]3'�ۚ�#*sZ�M�Ţ/��py�&��B�d1���v��XI���	���s�e{��zÍ��E� "��{��]���/c־9O)�F�?�*�"oDU!�)J��M�6���/CB<R\{8-��z-�TrrΏh���\�z�U!N|k�% �4��5N+HZ�J֕��
�6,�Ɯ���>	G�(o�+H1�����h��|䐽��F�/���k+۱�����0<���=�I)�?�P�䆿��ܹ~w}=�vn�C'�6Å�O�3.u�T*"�����������W�����a؏0�c�}?��sBd���)NF����Ns��MY��/TH�}"���"���ۦr"�ʁ��v	LX��n��(;���:7_�x�n�b�<	nEw�O>
lM�����mL�fE�&� T�� �3A*�ͬ2���,D�V�?���A(�4��G!�8@��0���{�6�*Yz��9
׭p�H`f��~��0�pm��&�P�b�f��crf,~h�v��j^_�� y9_��R���e����ik�5���\fӏgiz@c� ʿ��mQ�#�_��y�1b�i6B-)����J�C���νe�M韺.�/'+�W6�H ;hX$��dt�d�kr&���˨�����N����l��c����b[ꇆ8nE9���F�G�[]��I�)xcQ`�;_(��}������������_R7�������Y���k��Gdh��=YZhB"M�g��$�n��y�ό6���0��!qL�UA���Ԯ���q� Z#eN0��3�s��k�>��e��)���uO����������l aM�޵{��X=�^���C�#r7 W<h<m�r<��.�Y�Y<�]T����g.�*ⷩ2��Ȇ�ͱ5��Qڎ���+mHԤ	]Զ��$d�}�P������{�K�<�P��T1��q���K�v�p1�xʢR'E���X�
�Ġ�Z1�	������M[��J�P��8E��9�e�K1Q��t����Z��L�`��*�ƿ�{1h�	q���L��M0����Gcܚ�ƄR+�#��D[��f��m��"��"[F����#��n�K;�t�8�����M�d_��%����nu��G�5�r{Dm�E�z��bɨ���bm��4�=���� *�a0�/ ���;e���j4����/v_j(U+MC�n�3���^"m杽�߯�V�l��i��
aL9�Ţ��<�k�R������q���mUAZ!��R ��F�n"�:���Ң��M���F6�����CAbG�B�Ƚ���TU}5/�r�� Q]ɺ��G:ƾ�Ej�N#(y��I�P�-��|l1�g�o�U%�/��6�0Oׁ�0��<V
��1������!��9��j���>�9b�w���,���D�*�$��t�`�0,�m������QM���6�L��~��2�9:~a�[�AI,��=^�Pck�,ݞ�Z0`C���"�dm��N��}��!Yq/�	���n�L���r��I��;}�AX,x,�03&�/�ST�#pC常n��ά�� arK=�u�/١��5p:�Zo}4~]l&
�P�ܔj��ѫAAl�		o��E�z�I���2j`�g3a�:=$�(�C~I O�� ��I��)2�A�5�8��`�,���B�~x_ 5��WJIؽ�뙌͇kV�JH`\_�D���>p�@lB��� !�k$�h:��ˮ�৭�����̢gJ5 ��`�s���Gw�r˳4f�����Jgs:윕Q�ub����1��,p0E8�)l�� �]�w�{�ij�g�&=�:#�VsZ�Rn��jV6G�p(�N�!Bvm������y/�E�8�j�T��jru�ԩ?@�e>#/�FWB"�(W�;�I;�z^�Ne�|�*�)$���n�b����7&I����І}]�e��T�|ͮi�s�a#��$�y�۩�Sl�w/�yoQ�\����0&=�)Sf{��W��B1�С]̣�Z\�����rH�l�-s����>�Q^���Ȥ�&�K�BX�}�j��Hw���,�c���$+�@O�����'0"���
z��K��<���m����6ࡾ���R������������u�Q�5���fN!G�M�9ɳ�¨�Q�֞��Jf(;B#,7��`L^C�U����AgB% �~DyK�>g6!T�) �D�MK�%n�b5�9J�6��7�)���j�����4�OB9��� N�j�wS�4��*D�����٨�?P��nӃ�0aS�x
��Ώ|P��$ѭ�P㻵;|\(I`Z٘)�䓦�m�E�2	6*e�l7l�*��~�y(:��RMA�WG��vm���&��Y�`�����K�ɟ��Pp.!�,j=��<����61�<�Md��t�����=����iߥ�y�x,�lb�+B+����G�j��2L��)N�6s�9Y_�rɧ�?;�_�o��� ���+�q��rr|����+�g�d$��aiV��34��~S3"EBԖ��x��d�E�1
�5ǁ���j�~��(B9�7����!��?ˠ}\i���-Yx��7�.Y[oM��ˋh��(�k�t;�^�����rlU���.,��]!��=�ZyA
ig�c������E洳W���cbv��9k���>�<�N�m�8�ս�� X ��L�!��K��@ ��w��y��ĄJ:�-� �qUO��Ef������d,GE$=|Yւ,�)��{�����~Z>��Z$'f���I9lX"L��{X4	V��q��W:�4�qڷ�s�'�F�[�w�r��э�K�Xx+�x̨[&@JL��.Q� ���h�����'ur��/㵇��� !�qp���pi@�t�I�'����IX�)W���$K/ܝ=.@DS�{v��7��8z ��M_k�i�S�t�(�C6���		4��tr�|~@6��/��HR#&��w�+p����7d}��C$%d)E5����?2s[��ΧE��3���hϴ�1ֿ����o�Z��"rd<��z�Lbh�j =ª'���,C1���̓fv-�C �BN��8s��Au�Ğ�1�kӽ�������3�l�jn�
�} ��h�������O��/�'�HC�\��␶g��o�<@(ϊޙ�h;$�s�G&�#�;P4x5��?y�$&kT��D,!��Г��X�ʭ�W>�W��
���w��\h=�G�Ə .y_���q��%F��Lh��������������O�&�@t�/"���;u��r��sӏ���p%�#�蘴��C����p��-KX�ж������f���o�Cd%���|�P�!��jy��7є��k��R��9y�����,�OSᧃE�'�@?Fna�k�ca�q�vt�3��.�5�'�ׯ� �;�~�0�q�-d.6���#��r�T�@��kfŊ��Ac,�r�O�Z��.��F�y���(���AA/�>�P�Jo ��ŕr,����&��LzƯ���^��9���[d&�1�k�-�ې�a
�si��� [h�6XTY�|�W��ǅކ�~b�/�t��y;ߛ���I#QmL��W�$GZ�=Z�+��6���@��X�Uݫ_y�y�ɖ�d����b���X*K��<SRKם> �������o�9�o��{�{����9��1�w�M`��0�a1�̐ދCpas�Z�8I��vSCe�s��������]��4�q-��(����OF]�����v�<h�F*1�{mC�2eg�XXQu,	H.�47N��� %�{�!v
3��-�_ϛ����Ez��4+��nIuJ[��0���=q�ǲ�Uo�)�������ê���e�/��+B�T]� (����]�#L���l}8��f���9�um�����xZ�̦�J�ȵ�xMGt"<݊b��6�gx�N��K�J`o�nN���!k3M%y~x����{V[#kt��?���:ez�9߻�L�+ry燙&[��6�l>�7��9�sbx��P�3sX��[�5)[��O��"��N��I�l���]K� 5����ǉ�~t��!����h���B"NY<�I0�՗8hr�L�3�� ������4RJ�0#^�n�cU��)�r�����K�a9��KC�|��߃b���~�0�~ �$<�����,.j|�ku�u�����b�����}�<�ox��aDD9o�¾���X\�4������j��2V�G�?ߋuC
 
:�/_v����lQ��GS���z&$�Ԝ���X��>u�D��V�>0+�w2E�l�PG>��Orow���i��r���Г˘��Ψ~�O:�͑��j��	���^�7�?�K��%�Yi��ʶy�*�c/��{�qs	[N�JU,�����k&^�!�"�w��j�锫$G4%|��%fϥ�cU��iJh�E_@�W&oݡ61�� G����c�M����$'�#4r�@!��_0|^|��U�곾p�Qs�Y���Ū��ri��t���c�����4�XG���bx�N0G 9��}d��w��p�GW]ަ�/��I΀���{eߵ=k㡋R^<,�U?�p�b��
�{�0�����\g�:�W(��/|�	mN!��b��Q���O�Ha�3*Fƺ@��3���8��gğ�t&χ�Y"��xi@d:" J1�	����,��hAlV���tk�yI�m|�� �������f�V�rάT�UP�������ԩG��#H��
�䭋�A�.�(�B'v) �
�L�[�����z����:7�+\"�w-�K_z�H��RGr|YI�����}b����[�B�	F�t:Ci����S{1I2n$�J� �}G�5���׭��}�_:��9��QS�uH^�sAo��ڭ�
�8�ɿ�93_����,�dh��(�[��د��9�U�ۈ*��ɍ$~�CY���l#���D;����������IU�FY���f-VYp�pvP��cE	t1e��tf���v���Ͱ�NW� �(9b	��\�M�7�e�Q��ME�LL��	5��-  ��c�L�hnn�)v���������W��Qi&젽g_z%X��*pM��\18��׬u)�f�F�+��^`�Z4�Nk;�ho���$Ax����8�0���?��\��p5p��g���M�x�E���G%�
�O}�n�]�jG��y�E$�M	���t��Ǐ��v�j���Ud�8�D�-��|��p	z<|��w쎰�	�m��,�c/Q�H�H}�ҏ��Md :���[4C.r��������.t��P��&�Y~t8�%�7��>�X3�{���8�<po�_Rm�MҶL��$ԹC��4l�/>��~J�ԃsl� �~<��#׭؎�[�şp-5�D���� ����+�њ�n�pq|��X���B!\̳W�C��ѣ�-r?�dy�,���D�rEBI��]
�'�(4���^�����c
����E:`�i7�[e�C��E��6@>�5^�Xf��������|!�쒧?�Śl���I�$�og7dP�`�W"#�%��e��d����˰#G~[Lf�/�ͩ���>|>M�p�Jh�����"�x��߈W�����}�՜w�A1�:l��/���:����;O1�RI�!�u)���|Wx.�����⃨��k%8>��� Br������B�c����JY���KH����
�d�Ț��g���g�c��0-ۣ�F�>��R���T�9Ex���c��!p�!�`>�t@;��X�����t�$}��#�^R����l��*Y������mĲM���섇FL�pڞ�:�S�k��4'���$y�i��5n���y��I6��| ���}h4�����9�X�&;C��1t܎�����+�㐡��~���8��D���7�R ��:��[<�k�?��?��1X��}�sSe���u�Ϲ����BHW2|R��7���6I����c�a�q٤�Pi�嫋?�ծ&��$�]oY����l� ��0���+�~a:�edp����'�\��	�+5Z��5��X\L����`��S���%�|U<H�4�J��u	���q��� �\����aťl&(�|��\he4ڢ�����c��_<�P�q$-fX��GPg����/�A�WS�EF����1zy�/�;�>��)G�̭<蒔>�M�n��ƸN|U��G��uX l��YU�h Z������/�aJTMȃϋ�ꉻ���*Q�B*Uʰb7I{�)����R�~,�V!^g� ��a������dB$�g<'A���v:T#���ݲKB��4RD0B,�K�@�4��>�RAFD��W&�W����V�ZO���n�4��挓X,��˃e�����䖔K^B�JU�'�/\�؀yB���r��l�b��)�o�=zb�P�&�-�]e�1��!,�`�ʵ��'�f�"�ɓ"�t	^	#b��Gr�c�ʀMx����>�[9G^�g�?>��Gȏ��X�uXM&A������}*9 �G�G�Qd��-¼аǘ�� �&�;!j���Y�u���r|�����O}*�'"	S<��jq�#���L<Gldjy�1���N7 kp���x�uM���t�Ȁ[��!5���G����G�+����4E���K�#Цk~�i=�g1�fY��j���P^� �=�-g��y�</����D��J�½Po��[=�F3�#nE���;6GB�*៾-#x��
�T^2wg�<G%o�_�͜�l�oP�jB��hL�,f}���^�����6�����B����f�BV�12��.��m1	��t��8�d��}��&94M�5Ԇ,PhR��-JF�A���S�P�E�h-�����<��o�_9�S:�|���>��3��X�[K�R �I��O�by؂�e����W�5o�}��}�(�X�ҞU�7U�2�L����`�!h��AT���:�� 23�;��'5E���agÝS�U�O�H�Ռqwϩ��f	e>U��/����T���� N-��1���/���c�����v�J�F�DGtr,��L���S��L��W�'�e�<�>b��K��ݍ�s0�L���ɭ+���#��L4Ǹ���nCE�Ư!�%�V/k��o��:�
�l`�\����DH\F���]��Cx%�����l}���B|��!�ޯ�t����uJ��CL�Z������U�E��ܖ�jۈV�F1��Ұz�⧮�%ٳ,[wW�k%T02���N协� �������igѐ6ڦB�r�qX7��Fɍ_��-;S��}� gQL�O7��jj��r�'V�msVU�4u0,�8ۈH�'�um���J(A�G�m`�U��w��b���t,����zzb�3������3i/θ����H*K�M���F;��!��O�)T���q�kۮkf��uܹ���f��c����P��g�� �"-F��zo������<L��V�%+��Ģ��" ��&*��s��I�AB$7�#���R�����} f�?�w�'>cƪwnrK�����(��.�52��+�7K�U(����8���ێ?��fwD�3c�Q*v�j�����|Pq�P��W,H.3C"�`�	��v��������
yݪ;�η��u�ӳ�pb�r�C:�}@��Xo���\����0YN</��<��d�,ov��Q����b�[���v`}g'�d� �d�YERB�U�����xF�"��1%%��gf�[��/s2�t�O��i����T~�Ra^���3��g����[��c��PU�,�<�F�2x���r��hX��u�Z2.�\.���6ea����:Ʀ"����[ "O��8���Nv �5�f���6*�i���oy[��\<�����{�Y��!wF�s�����GT���/��@�����d�LW&L�h�����Jj��J�`��z!7{9��%�Z��`�]���khb+��2.��qP�N�As�\�Rҟ}�
��!7�F�L��t��K,9�=���ЭHv��U�δ��h�'RU�,lI%�//C�!��K*=r��`����bD����� ��1���O�
	�8c}�]��4Ik��-`]�d8HP�C�xZ��.����$g1ʂ�&R����Om�R4��ZZH�(N��qO�r���t���<�Eđ��f�ʽ���k�����#I|�2�R�m����&'�c)���=l"�+w�3�nu�6�=�w�
���╎{nm�R���9+�����"�β>�}���[�b0+���Gt��rYxI��g`% Lv�Y�M�].�D������ء�wڏ�n	L)xUުG1} j́��ӓ��E�^�]�'�������U<7%YK�K����԰�-�v��CI��E��"���ETEר@`�(�ɐ�V�&��D��o��\����k�)��IM.p<��|z-@>P�c�d"g?w'�e�ٷ>8�S���p�WFT�*�n^e�P`T��H�����WM��d$�`T`�`����+G��<�[����̦i!��p)��1\�|����
�7+'q�Ob�o�hg�jW�f�לը�o�Fq�&�Y��Ј�G���.���V��yF8\�e���6i�Þ��tW�2���^��!�b4��x�OM��/z�7�zC=x���&��u�A�8#B�v�H�Uw&��Q)V�Kx��ݓYo	ʝ�m;=G�IiH����7f��eD	Ww�]�3��U�a�6R2�1<�ˢ���==$w�k�8���������~���;Ә�tn���au�=i�-��uTv��9x�P>0������_Y��Й��r�h�
Ij�/;�6�Bz��:j���Q<�	,Xdls�9߽�U��U
 c��K���f@��4�i���)�~bǯ�¾�>� %����Ym�{�*�qoY��p�Y��1ܬ$
�!�A�V�@�U#x��Y�6#|�j��R( �#�y��l�ׄ�U�z}�H�@5����Ԏm
e��l�I�A������4u�x��-��`˯>'�]g���SRB��T=}��]�IY���7�_��H�D)'V_���؋����A	��_˛�#$�x�ք�z�
��Y�d�K�D8z	����+�yϴĀ����n�qs��q>�D�v�ͯ����W	Z��7�2��z-��Q'J�(O,�Vȋ��+�m�0�V�ޮ�U6��USᆳ�"-����>J��#T��)�
qt�D�=-�[+�3 ƍTVE����B�XK��;2μ�|sr��\O��[�9����_B@ӭW��1h�_2���{�rq�#ſ�M�%�_�F�R��K����� �� �_n(�̗;K�b��8t��%�G��+Z��œ����V�V<)�-���_y#����~~���[ۮE��_�	���+l@υ�-d&*S/��|V꣩>i��w�+�r��>��v�s_̳���?�4��'S4�*6d��1.>R�^��i��X�je�K@�=�ֱ���z��P̙�f����G�٫_����z� j۪��4@Bϓe�k3k�C�k��������2�����	���~o6_Bӏ��6'��K�E�c�G�M�u\8�7�D�l�Dzi�O���R*���#�<��C.�s,�����R�`b%�KX�"��ɜ�k:a�^ĸ��^����l��2���W-).Q�����V�6+�Nl��"<��v^��0�̒4~�4���)@MI��uP�VM�Ʊ,��~��X��NV!G��P&=�.#�� ����7GQ��etAq&�1	�D��*��kDY>�z|�b�<��!��D��oYE7jAX��֜������qN�2�<��X87=O'@of[6Ӌ̮�a��h^OO�Pw0I��A΃�����w��C�wx`ꠌ��׺���V+@^s�y�l(���J-�Ѩ�ُ�@P�n��ĔP
o�/�i�/�oRH	��.ŉ�Ӓma2B�'�F����]�(J:�����������%��F�c0OI���@R8\ 9=�h�许m~cq�jA]V���PqFZ��u�X�=+�X;����T�F<����£�A̝$������#Z���8���C���j2�*�r��0Ùѯ�.��<W��@�'����m��z.�}�ՕPQs#���'�8���L6D��>�ܘDX ��p=*� 4ҝ�V�.!��+��2w.`g�4Y�:E�A��N|h]z�)�e��8���l�OC�Ե�-��n�s�IS +�+��-�IYb}������Th����Ȧ����4`���sh'UϺA�
�>���hZ��P������w-y�S�Y�d@m�^��5�}Pi	ܝ���[�q�VPlǗ�p��ȌlaR��_�6��Z׊�n:�C�M��ޔ��#\�{��x+�^23�T���KA�ʤC�yقgt�5Mq�����^!e;yܜ˳�7�~0ׯ9[���a��̐�cRTO�!�e�Zs�G�o�[0|�h9J��X���ʟ�^w�/-�MB�[^)�)A�TK�O_K���m��x��F�0��!5�|Ėf^�B�`E[�s3��{��H%�w����3܀��8�G��:I�ay��B�sL���n]{�|n�e�|����Ԙ�jU���Եud�X�T(��QX5-��;����-"��{��UV�n�)�2$�j��ҧ:冯O��*5Ȟ�Cex6�R&�q��3Q��~g���5�:E��8��)�p�hxz��(�Xx��c7�F?Y�ȡ�ե��M'e��UjMo�;6:-'��&<,��Լ�>oJi��,M�$���<��F�y���̯����srBy����W�O�� �Tq�y�j��9ǚ�3=�BD��Q��I�*I��|m ��g�3���ZSӖ��6��W�&��V7�6������Ig� �׆]G�y9"_C�������y��GG��«	I,,TN�L�wV�yd��$�~��㡆�ﭦ��h�o���=��Mo`NO����7��a=;��A�>�3�0+
�Nn���3QV�g�2`ׁ�� n��/�~|VXA������y n�x���B�̄m߰�ګ��DH[-g�ۅ[|l�6�s�)����r����ҳ%9����sqoʏ�`��	#��(Q�y�� �/��U�h�r�(�UUyp"Y�$ׇa�bk���^���[�n��3-���>'n<ng�����Qc´=�Ѱ�]�'a�3�a`~7��S�,�:ipWR�7�Z�L���u���ں3��;��P�_hpa�x���j�kq~�$>��m����'����eӊ�sYj�v
�Q�
������B����I
o��Z�ך��[��׽�9 ����G`d��%5��?�j	�EZ�#�� ����c��`��r�)������$]"yw��|BxW��Ӹ��v�GUmb�U%��_Ӡ��q
�-��s`=��+P^�5}�<�h	�$ݸ�wF-����jO~�L�U�JI�����A^s�1R�������J2qd>�Z��?C��`�k.�v�FEo�� �qZVtd:���[�y��@}o�Ӽ�z��C�v�1����v��^�[��/$���&�5��樃6�9����$�f��Ȳ��.��@"�b뻼m�Y�u��`a��kQ�.�	}��"��@�]��oKO�=^����goJk+�-~,��<۹�p�h�QF�4Z,���D���N�A;��Y�t���#�~wˌ��h������8�wȤ�(^���!�s�;�A��w��!�Ƶ�U/:#D����7�����M�Ht~/�tB����=K��T���rZFs��/�h6�8��`OE�o���vW����T�=NQ�c*��C��*�5�)��`�-(�T�M�nD2(�����O�Q���
�q����E�1�5�����C9� �ex+��	kaKl��])��춝jEe�����+o\��EBm�F73�����:P�*r��g>į#���Fӄ�4�� >[�Пj���6u�Sb"ԛg�f�jT#�B�(W����5W_��x5�~�h♪�Si��[ RΘ�,�F�! Ӽr�I�
�2���p�ko�.G�5� ���ڄk�x.\;�f�/k�<��8)�<+���ԀY�Z�p��*Q�_35z�}����h�O��>��e*��FM��g��:����؈�R�l<d����C�~/�T���=� ��zs>�Fd���L4����V us�I�22����O�w��ʡ`W���H+��4���������q�u��́ �sH4Q�e{��v��տM��9��J�h�ើW~PQ��h��С���)+�zs�w#o/e�#�G�����P
鏢P53���S!1��z�rN�q��C�lJT��} z�L8ʢ��|�M�+�aՈ[
���M<
�����abɭ#�N���;��?-�cj��l䐭�o��k=?�!�.Q�N�{?IR��L5���N3Ǥ��.5��vM���e��-�z��8O\�6�ԝ�[ʨm�J�2�q����4^�߷/����F���ڹX�3{z0`Ɍ>��F��9�L��#Yt��o/d|�*����A���zv|FqϮ��9w�8�v<q+'��h����INs���qB��r�}<��gR0��[�D\�+����pe>f>2����V$��'<gY���ӻ�8�Ջ]mctd�8_#�M�������	l��m��0�]��k(���t,dO�`Yz3d��QO-E蹒��b�vW4{ּ/葳�kTK@Y�HN	��g�v�w�<��d+F��R$e�	�tR�>��xd"��a[��2��ؚCQQ�o�֡mV�b:9���	���iu���	��&B��L!�4Zq��B7�g��YMۥ�{��}CbW�^��/��M%�'s���T������F�-�{�M(����p�0/�.q��:���>��^���.(^R���3��0�V���m��S������aA)���@�XVK��
m�3K��8
1�#W.�$U�Bs���+S2���z,6j�$��2�P�qT���S�<?��`a��� _Dݟ;3�cR>/��V��d�͚L�hХc��	�z�գ��X�[Q�lB���E5�y!t�Y5�#�r��9�IeYV��,��7K�֩hd���;����,ί��<��PP�����T��z�eg½+|���p�L�J�����BL�i����a�p�<G�y���St�g͘No�o�D܇�9��h���D��Aq!8��Ur�%=-�d�u;i�S���!~x��$Yf���K��-�����T��JB��|0�!Q-�qZ�'��(`l�[���Zs�oeu:��~�G�~vKp,���3ܽ���H����{�ݓ�J�/�0v����U�p��j⃥RmM�^��q敂xЭ�@���ı�r��p�\��{��x�b�D�E��inXｎ�f��f�^hc���T��ʫI�\0\�s�A�lu�t�o7�i؜�3�~@�欆�~���T)Oa��j�aJf`+>�ŤT	&���x�;����
~t����Z�ޢB�z�L�t�ku������1���}�"�|k�V���:MB%fk�ge���P5�D\��S䆞��&���,-l?.��
�E����C��>�+�o�k��G�FZ ��yN#gU�� ��� .��9U�\��D�j��p�*������2,�ѯF� }@	+E�O(5�6�ҹ��ގ����izhjy1ѝ>j�b��|a���q/�+FT��9W���V�4T/�&�_nŶw�M�k#^M�MLg�-�Ht�tW^��qS� �A���F����f�p�$hf�D2�"�z]/dnK4~ہf��|��8��O��ʿ��d�1����ǳEb����L*�&��P��	�CT�
9�7E��8��kҔ�(�":��r]&D��޾?]�J���B<� ��Ć��>�S��|�Ӆݴs���(��L�)[U��)��U2)��ʠ׻ǅv�i��@��NT�������͖�*V������H堡yU(�xЛ���/>hT��_�!O^��k5;+�Nf-H��ş$�cnv��z��5��.2��g%;s�yb`w�R�����&؅O&�x��k%G�@N��;:�
��8�0|��;^�|%Y>�R^�H��V%9��M>O�"L�)s���y���iN��
��O��q5�I.b~Y�:7�#�8�)��K�5��N���1Ѵ���P�D�;�'��\dH9�g�'�lw�e�Bx*2�5%�R�0�=H6�-Y�����������t�An�W���%�T�4@����_Bm^��)�)���FR� ��6Ny�"����(���f��8�_\N~%V>��TZ+'T�qJ��v|��#��I��2�?f	��=����kS�o���X�,�S����}�"3��|1.l��V9׋1�*��I#�ȿ�ӈ:�$8P�*'ļ�t�Y�q�k\�
P�3�C����g��\���Q�UV���?�N!�8 �$��=S1"A|�B��An�5�9��0)\5rJG�����^�zw���D�f=�W(	�L��<kr�*�H��G�mr~� ��"kJ׵D��9>,���Z��а�%b۠��EɁ-�j�
��ɇ}�Y}7d��KHn� �r(gC� �����@)�� �I^�0OF�}�$�K��f��WG�x6^/���J�';���br��C=���ɜ���(r?y��lV��K��w�u��Otdv�rPK���؂Bu�Ƥ!���B�A�t�h���T��`��d���V�^��z���3@3�;>*�%�]�xa0��!�����I^o4A�:�pܬ��g������r�@BE��/ɨh�$*�<�H�T41is������X�7�{`[����~���!�]-������#�h�=�x�&*����p�`I��`�Ž��F[�*�P!!S��,�S��7��*����P��̏��<M�*�w��̠!Ó�o����:�\0�+^6ۏ�.5j�0��f�#��B�c�9�̌�2��z�E�D�Ou���2:X^���g���.��1��rr��`�����6ѕ��E��pJ��#D�:�B���5�m/<ζ����D[)�n9Ut[���NY���k�6r?jvj�Q'�#�i�����MB�Ｒ���]hS��<G2��M.M���5&��5���:rV� ��'�9pD=����PI���W#�>>� WVRC�o�T��X��ޘ#���.�o���3	t���:�T�3I}h���],l� ��}:���XD9Ȋ�B���<���Q���w��s���{)�گ7<2��6B,����9�
2 &���-�j�J��N�C�]
r��as,)Ռc�ߏPU�v��������?���ۇ=�	m�3���eO
"%gG{>�S��� �'�m����aoҙ���Y!�ҙ��	�p~rUЄ;t��

)�o�mᭂ!p �z��N�%� 1�˒-�od_��<�c+p[G�"~�R|�@�z
'l�14*���['peĞN6'#��Ɯȇ]sx]&���m��B[�x<���M���ਕ�Ew��#,_N��[��H�-������Byʅ��weQ̚H�����K xj0�g�J�J'��朅��s����_�(������ 4��+Ȓ���,�*Ts�oQG���r�WC�q�+��D;RrL����.�#:��� �!+�PIڍ,��L�����T��*����^�czǰP�݈H�9�`hGR�YR�x[�:��y�-�"<-?!l���!UBXK��;��A�d���z��O����8��@�΄uy��_W-���	��*ң``�P ��aN���ӉO��E�&�Y��w]�I�;^$��W���x��U!�>����[����<��}�)te�;ʴr>�?I��#aΑ�uJ)z�)Ւ�����6T=�\��j̓��x���ϫ�`��j�=���s�М
İ(`b�����^�Mc��vz��;����0g��S4�x��M� 0+�`�����T��3m��\;O*�4uE�{����P럢��<�Ci�XYs��x��\�:�ܖ1�X����Ͱ�,�=��rr�l{�8��ܨl2�����?�(��%�H��u�{صc�$خN��-J�?���ם�-B%W��,��ԼjCL�\W~X�{�U�o"�/jLH�i22���YP]�M���X�'���YV�
�n�T���'�� ��9�����S�v-��H)�i%�Ȑ,�",x�~�>�/E��7��/��O���-����I�!�`�%���w��f�0[��4�r�o7��}�kd�
�7�S�H#`���g-.$�x�ϊ��:�����j@&�#���[��&��^�\�������S�`��E��C�5���G��P�;�1Z �2�À�xkd޸.Xc}�ÔCa�ڵ��Ƕ~�'�;w�T��l��-�ඁ����ucf���&�oK1�`xnY$^bRb2��u�x�۝�'=�B��
W�ʫAs�ƻ����=qPB���f��w*�*��bW���p儽M��4�\o�0a�>w	pF�2с��!L4i�����z;�Oa隷�1���Q�=�V���$y__��s�Y���{X�+	K��k�cޮ�`��޾�(�����2�҉q�������v#D�gA��*��;��6D�r&�����㦯Pk�.h�~�(��R5�Z���������/��֗��+�ooj�X5b)U�p��v�3�}RϺ�����^���@��
���_(X�j��20�/&�ŏ��9I8�Q��E�[MS�����-׍�]qX��&,'�0�p&�'L����U�w�j�D�c�Q���L��>��\jS�Jl?�*�SD:W�Li�7�TN���f����f�z���, �b��Z�=�#���3dU�5`zeW/+fM�b��ɭ	�LB��dÉn�]}��~<:��޴\?r=�&�N;NA�=����u~��rc�0��z�i��0�ؽ���q�JM�V��o�<�}.�L`���ɒp�	;C�܁v�}�x 庑i\!��aiJi4Lt�O�ϧ��^K���OB/��: K��]p�\����e?VnOD���ɟPFJ����,P+@�l����S�Cvq4�	S%��M��a(:v��[�l.�KB)X%\�� nN�mq��V�&=����?�h�x|a�b`�7�x�z�@���e*�~����k������y��w�)��wZ�%�7�/P�
�<�A�wC.ǇF|,_��x�h��p��_d����7][����E��_ݾ����3�� �{Gt��a��F"�wX?�,�����U�{M��#a�G�����TJ#��㕁o�T�Eny�6��h)��!^�ڞ�8` �4a`���`�c���8�V�x�@oM��Z��? 3�1�w��%�oďЗs�����O,F  &<npb����ҋ ��A�^f�3nE愾�\��h����f�2��]5��`	��2���
Ҟf@:~z���W���3s�G�4A:C;�;ߌs�`C�jy�����rY�p�VMB��ʞ��;�B8��ˁ�ەq�7�A��uy��4� �&l�+c*�|��A�G�4T�^�0�������	o�4J*m���ۋ�2�w�<C�٢uq���'u��`,��MA�b������>3�Iꕬ�4�H���8�)a�x$���^�ܱ�@:�\�HnO#�?�'�f`���G��Z��"����B�J��"��Q�|�q�����o�Oђt�V48�z$?�b [j��i�Һܐ�1G��K�]:��O�4�4qqN�_��,1mg��v]�6�XW6�ꑩtC9o����q=k��}Jx1��A(���oKaL�2��_���!� +������NH��IF�3.��uZ�a���#��/�g��}s�q?n��SG����6�N�T�~*��GK�k���5���~x�W�!挟��B!vFuN|i3_���F.ߝm�O��G'?:o�eϓS�5�cq?�=�{���(N�5�O�蟟Q��������T���k4U	`��F�i��[������3��к9�t�UΈ��T����>�w�� ����S$��U�?��vi�#��3ޮ��u'zm�lT���d!h�(+ci�����!Կ��:�۾�JP�f6694�C&��&[�=q�Kg/�]$?m�+;T�/x�ǞNr=�
.
��n�tϣ�G�b��i:W!��D�`W�9��v��_v�O�ms3�50�d�B�i��f�?V�*]��z�Aﳟ!��s���.���viIU�'Ւ0R�\J�sG�
���������״�B�,h]�1d�n��X�zs&�3S5�������d�Y4�9�+�9Z�'_�z�::6��c�T�p�`v�<h*&t<�A��]�=�Y6�;��f�$�"sԏ��GM�[���rt"X��ٚi��S#�+��m�$=g�7m���k:���o������>n���~���# ���5ؔ_��(aWlAS��'�ǡ�ܽ^��T,��Q���IϞg�c(�-�׌�>)�� �1��cy�"m���~�9Up�%�?*�x�,��;uף"&�CV��X��F���(�i���$�#J��0�W�R�.��2���Y���S��~f����ޙ
�Y����?ypPґA��0\ܳ�/lN;�"�5�^#t�FPE%�����y����M�|�"f���vpi�/�1�t�Q�aZțe'�T��ׇ����QB̉'�;*nH7��;��������񄱋��J-jn�p�IU�;&*����v����C+Fܶ��r|>O��E6�ie��d�v�֩����RI9��.�R�;���7Q�s�qK:]KX�s�I]��sQ�޴�*9F�Hא7�-ou�vaI���c6U�������áz/m�ܢ��؅�g?�{`VA��sg���߇��A��b֬!�(2�y���ո�aU6+����+�P�����S��F�a�D��d,�������܇�D�Q��a���<��!��uT����2�yJ�����O�·�H�W��:sDځ/M+��b��SP[4���2-q:�%*�� �b��@�б|���@
h����Elƪ���G֑Z1z`"t�&����X;<q>�A(\x1�����C�c�"U�\�ܢ��8#�������XL�Cd}��GyY���������v�O�k*��%�y҈�?(�������4br�Y�@̕��L��VJ餽���qk�+\��z�=ft3������C\FU��r^`T�̀�4������
YM=.�+R��$��%�־S��
R��J��S}����G@��A�T}���❅]�~�?˺�8_!,�i,�~� �Sm�f�22ަY��+��!gLoT�m���P�~o�-�{�d9I�JU�����RBT5��oTJ�|���|�:&T�C�P��>~�N__b��ѫ%�3����g�
{F�����"v��ż1���N�lPz,-�Ҍ�����Ղ
z]$l�T4g����H���zkX-J����]E҅�1/��9oa��xD`��P_j��F�t��X����&��\��������3�J;,rQ����\��-Ja�fF
�y��k�n��-j��	���G��&����y.�eݵ�Hy�:C]�{�E��vÒ�U��>�(�M�#q1�0ʤ[U�'=;��E�'-��f���"3���U�ຉ�+�$C���ϛEjY�ػ\���հ��|9;T�7�_��\��릾�F��
x��.�*F%�ߝ�����ui-�P����|��A?{Xh�����f^��X�|�s��Dx"��R/���{� ���ܖ��h����<Z��F��
$���g�Ώ��"���/��ߍ�fff�1C&��'�2��]��FYn((]zaU穅N������ڱJ?ay���kB�BsK�?8�5���G�]��#��z��w�a(dKf7��jp��=�6�M��}�4I�J��*G��Y�O�{|�*�����d\��J�	�Z����ꜥ�����ȟ��F_��4�T鎒M˃�HW�!��,5��aprB��9�߫h՞^�q�%A�F���r���]�, �h�\AF?��#]0���;��Q���F���K|��v��fX�Z�����*n�jt�^hŰ>ϖ5�:�uAIAK;���R#Ό�6���K�;�u�t��Қ�"��;���VL����QJg���vɌ�"J"��K!K��!�њ9f����;�9,���0���W�H���k�����S���ҸH��Q�������wi���ft�^����`�W�LB��<��=<��;0)��@ڭr�~�������bl�Y2��~�n����J�u��Uû1��i~������is��
���ZPD�V�;|���������2��"u��x�F�*]��S��S�J�F�K=���Ԍ�)=�*�`�?&7r���9&�z�k��?i_��'�48櫶(b�� }���PrF+E�qT�s�OS��nb��8��
KPs�/+/��nߥ�J� nJ�/&�W' ~���$��x��q��|������a�̚/P����sR��J����R�@T���d�9ZӃL�hG�|<I9��k�yW�����|��H�J- Œ@�J)r��LV��3t�\Vo9�.P�`^G��y�|��B�;~W��m2 �)~@|,�w͛�8�b��f���P����ÓkJ�D,9hF�}X�|D��1�o�9S�c�Q��f����_��"�t�ഒ�����s����^ �a��Լ�s�~*��*�y�e5Y��RZ���˛�f�/�>�h0L�-��ugs�U�f�(,L焽���6pw�ro,絔�- U�[.�VFl%.B��&�{��p���:{=��5/��G	��֎���aT�2�+I[$8a����,`A�ɨ�l���%��Q��?͚�φp��t�Q�,�640�QN(�\��X�j%��B�3VsE�gX.�Nt.(�w�2i��"z�+WUY�T^���_;��_�=�g 2���+�`�='�bE��9p���9����s`X[|0���B?-�7�_7kp��L�2�%g��/: �����$>��@O!�X��Ӂ(�l�ñJ*d�� \f�'��x��?L�}��v�0���s(�W9?�5
a��L;���K�X	g�ğG������~n��66�@f3X�Io�NBD��I��GR�����舍傛�ث�JJ�J��k�f�r3lS��<�����v������J̔�4�߬�q�Ҵ�b��:*�m�2 Rl-VI���S/���������[Q��/�pʡ�Y�m��|wZ�Xv�	sA�b�]�������y����� T���%㤙@�p���9bE���b�^\����V�G��G�z��c�v]�c x���#\�Roίߐ��C�U��m��@m���ԁg�u/ � ���x��_ȾϚ�V:�ԙ8仿��7�MAWFln}�ˡN���
G�?:pZz}_�M�+��z� �V�� �^R���Ґ��N�r��S��F���ؘ��q����$��+�ႝ|CJ���f�ۏ׳��x���|t�s�O�����������lnT;�B���d���5���qm�տ�n�2�hIR5�_G&�J$�dΉ��d�����3���Ze$�ո��Ð���Ĺ�};&�"��q��������U&5��6K����{z9�Y��.Z��Ԅ��[:�"V�l'afz"u�O�DoNP���RX�v���hY�+Ń��|Y$�h�y��f	��c��t�Ck5�F�^`��$�2x�D�Rݩș�>���ΐ��L��a%����<j���""m�/eS(������/�	���4�d=�����z��;?ݬ\kb�����A��^�n��t�L�Ͽ��ֆ"�~�A����}�G��Sv%K��`i���эj8g_�R��K�&9�"�n�Ɣ�-\����� �UQ7]�o�m!߅������y�����������?S${����g1;Aۼa�K���s�� ɀPJ��Vq}2�)�WR��M[���� �쯑o��o�6�����;K��?� �D	�k`�I��	��9���7�$D��\����b|� ����|j~�=0F��@)0-�`����Ԇmx�C[�$@N����Z5#���������sH�s(��e������M|d�[Tт��~�hfjlU��ޟ?y��6I�ՊYs��!��M`�M�mCU=v��=��<�����y��;��VOC~PHI���cy��Q���R�����?�o/��E���?�� li'gM�촀#4�iVD�U/�Ff�T����{�����ǂYy���|ʹ'-�u��[���u����g�_5�Up˺�w�� �Rk�/�d�|���a����L�ܡ��}>�/S���O�x��	�V!8d��X]3YS�t��ݒ�	����oZ���(��y�K��-��/�^�a�O*�T��!���^���,4T��{��(�`lm�ވA"�I��
j�ĒӐ*�ܻ0
��DKz��
J����z-��*G�r�5E{""�C����c����Ğ�`k:�!����Įg�H���IPd.��}����"�מA��a§��stShQ@��Y�i����zC�
x�غ��eߓ�Ծ�ׇ��·���0�/�<��(��r����倌�M���u5���ܒ0��^Q���1��Poټnϒ�B{��͹��8�<��:&�k0<���-ߙ} �2�f�O։V;ݥp�؛��h����Qh[|"��e��~8G�׈v�_����I*A�r�t[x��_�R����&���Y��9��w�C�ãôUdI�h����^�^5,<a	�G�7���#�� r��,ȠGx�K[=�D��'S^�_��0�X���3=��W(#�{$B�Yn" ؋�v�.��oQ_9g�)%`SI�=����a�l�]��+�ۇ������4Jn+�cȊ;_:f�'��e"��ˠX� �>>s��Ax���;�i�u�e�zDngzY���S�<�]�%|� Ԋt���b8��^�ջA�J�bq��l��N�\�������i���=4��ݾ�k��I��w ms��3��g }�v.d�1��gB�1�����
 ��0����{���K����%���Ǿk٨4j�Ʊ�6���_�K6��M�������i��Mrm���g��x3�	�>I.�:Q��F�x�R��  d��UosZ7�r�@��A����v�q�7��T}��:�mx����T}�o�:�O!2TH6(AQ����ϛ!�����=�WG��ŇHqu168_�99]����T�d�\�ni�������
���H�H��}g�Pۂ�⺬�#E�b�F�Y�0а��n�'���{��������49�%hh��VАD�l����x=Кe�D��L@F����b�U� �kIR�Q�I�w��ԭL`h�n�Q/�̽�!*�r-�x.d�Ւ�G��C|/��/���:��ʌ����襓"��J/!�A�8�PS[���7!����=�K�~��9�,�@�p���ƚ/^�ot�ŘL0/G?��ك�nAS��;�G�=�"D���|;qgn��}7i���x�X�촷�Gr���zVE�-�e>C��6�&	�Q���$+���w]k�µ��b�K�ZU��c�k�a�<����s�Z6��>F(���[�??E���mc���@���Jg�G1E����"��3�/��鹩�E�OP�d�5�*;O��f�#��-��c�OYְ+������n������Z�A�Œ��+籗T{�[@����3��v�0�ԙm�^c_�+�D�`��VZ돦(O�O�~-%�#2���U�8?�?�k>({v�⛡�8�DOx?#{���J���o��R��h�g���dBh���BT�����Ǒf��G?s)AI��a����;��=���[�vUvn�F��c����ȿ�y��hL�{d�$Փ�-�~3�5�Q�_���Bwd,n���#w!���y~z�!ojJл�GG�1�!1�&i���xOxy}K5bc�n"(>놺�2�9�xHN�2��-��7�_�+g]5���KN����[�&�s����kB��Q����� �����5뉣v@ź�����o?�_&&i�\^�s���@�H�R6������j�6�W�׸ً3�Ƭ�.���q��vI"�6��fA�A���<��(7H�2aw����nv]���^��+�+��V2�6in�<�>"iJ�uu��)Sv)���{�b��=��i5�\WX�ǥ��ަ�2ሇ&N&�N�<B%�֍K�O���TR!�2;�����9�>����PwI#�䯊Nf�d%p�]�=�j-^�-	*S��K�c���U�U�,Z�o�}/��o����\��[��!��,���g %8�D�;���!Y`��Uu�Ue��si̳J�n}̭����@J��C����K
^}8f갿#3(˩����k�URx��@6u��HBU_Pm�QI�NE%�e�)P,E+�Tx�mO���P �R��-Y��J="�˱�`��DR;�E�����1��L\�^WV�d}��f���vq���:c��܃K�$�f\+Z
E�ZnK��s� Z�Ԅ8��F8�`�(�\s����Ҡa6����m1M��e@S�YSH7�[�:����]vE'��A����*[��u�!�T!��9��g���z������H�"aA����w:-�5+���z.Ԭ�� ]o���6�'T��d�<�hpz��S��HCv.�Ґzn�+޽�9�R�>�9mn1�`��
�;�	d�Hn���R�"����`K�Z#/�a��8C�v�Ear�#=+�$��inmZ��H���˳���k[A��vݗ;H~o$�����Ճ�#޶��F�'�����O&���:�zf�HLӀv��ףz��^:��$��My��>}��ք����=��f�_?�����֘����9�3:���B,�e���7�@n%%*�iv�R�;Yd^mw��_�w���sa�v������� �	�uR�3,d�r��_{�>��\�4'?�Hݕ6D2�s�E��o�+^}���Cا�rK��t넅J\d7�ح�uЏ��@8�O�*�æ��s��[�����:�jI#�os+��I�^^c���o�R������0q�_��1�e#���,�����Ӭ��#H~˧^Үo���&�3���f��s��㦰2�?A�dT��\u��^��#� H&_��J��rsx�*���տt��C�:�#{�L����M� �.{��G6[X�-��~���>x.�@카k����� ����(Nn*�+'h_�b�BVy"E2nTuj^�5<�B��V�mA���`���SHr���|��%��0Ye����px�W<� s9�o�f�`�n]K�c$(�t�g�?�X��֑�ЀX�Qa��jc[�]���*��,jxo�&�S���V��
;�l��Fȿ0� �`�dm-�������X�w��Nˤ*5��9��!���,�2* zLIU졥�Y��� �h!9/�1~��=4�ёe4�K\Sp;���c�r��GW�5T��=����7��EVe�F�Z���x\�)��_�'Ɗ���
_���]��H9�RMU�L�ނ�������B_\�jkxC���I��3R�ƥt>�}1g�-CLB�Q_��� X�H�=�t��<(l܅��JPL�	c���Qf�s�����^1E��(��<� CB��'r�2��������0���,6D\�?�z�73cD5%Z,��%�'��6a/ ��Z��')�.R.j��ol )V�jȣk��
k�U���M�[o�#���}�W��,�Co�({l�c��@�:��	@�w��+td��_Ф�ڀ��'�j��TT�;�	׆����\�ՠ@E�g	?��O�^J��I����:uqp\�q
F,�-�%�J��j�qZ���9j@ž[Z3�u|:~d�q}IP��ԣ���@>I�'P��"�t�Q���3A���~mb��)=���-�l�������hl�oJ!��!���I(2%�+0K�c��XGj�yx�,i���g��/f�"l���X��⟐�U����e�`��iw�G�C���J#��'�H�W�0����Q�fu����&*��H
 )~��P��Yb��\J�dR��5�����jK��N)�+� }x���ώ�h9\K�:�EJt�1�O<fLq*w�rr�-�͈#�}��X}��_f�ƛ\:ʇ��;���pJ��=�<�B��]qpT�wKJ��B܏��*�d9�R��U��$(.��I�]>�o��0C���x4ݼJ9�3Jd�$0*S�,\��@��<�~�Eǎ'�o�kљ���w�<y�������>�e��_s]S;Zfj��<Jh"�1�_+w�M_�V���3�?��✕��bJ�Mإ�mv{��r�w���#</-��Gn��^�p�de7?/[LAi�w��|�V1G��Ns���g{�	 ���/E}��q{ s�,�S	�hu�9C���o# ^�w��^xn����P5�R�壺�y��U�d�a��W�V�|�%$��^��Qb��j�1V�G���i��j(�N��d]`��m0�"��������X����%��}�Š�<�7]��뇭��quI���9%1��eJ����5�mCmHB	P�h�D�YC0�ro�\q���Twi�3�J|���5(��9�1���QJ����V���ǹ ����?�i�XWZ�����sެ�����f%��L���ؒб9hG}�}ߤ%nF�����1������q�0>�� ���K�z%�Y�YN�@/j-����8S�O()\�i�7���s�k��!&�+�U�G�jҜ}l�^���_��"���Rّɷ�Ϫ�������V��j0��&xH�iH����b���X�\i�۬R�M%��Ǜ��I�|�����[mh�]E-�x�bЉ�A��\�$d��ݖ�'�""<�������A/M:g�����z�7�X�r�O8���jC�s�.�A�!��;�^�_�pW�~�����]�����(�u-�V(��GDv����pX�_���������j
z��Y��-�tn�1"��.?���"�$�	�͛pg���܁'"
C@,D(e�m�%y�o\nK�a�*�@7��([sN���N�
Id�1u'Ͼ0\���h �m>� �vn!��-ᤢ�,a�d�I���+��Ǟun�	7�w�ϓ�P�|i�sFt9z��
u�Um3\���Z ��i��l�ʇ���K��ib0M.�}��m8��ͳ�CxIx������O��q�<W�LA����}=��?�����챌)�d6�q(��=z���zdFvʯ	r��"zvƅ=��n0<RP
L~���{�!@��m�\��'?n�p�wt86IZj��c[�{�q���É��0�H��}�m*M����]GL�x�Ж��*\�r�l�,2���%���>,��Й��s�d��Ӿ i2ʦ��M�#DD�������i%.noR4W���"i���m_��p�N7O���qчR-�ln�O�����s7� ��cXh�B�B��TC0����+>��mп��Q�Kk�"f-���jÊ�;�"�b�ڻ�m�����D�p$������أB���G�!qc�Fl�������n�P�h/��f�O?�%��H;I�d*WKab@	���j~��Ym}��{@L�=�s�D�7�� *�|I=
3�5�w�㲝� ]=�=��cs������V��^���?h��TV���� a ��p%ܐ~U43�}VJKe�ODR�cc�%uR��/���e�c�j(T�|CB�N+6ƕ'q�n��k�'�H��
HcO�&{��T��՗o/����Ty�:���ܜE�������E?�ٿv��5B�|'��E����]����p��d��(������wA9U[��ڹ��x@i�8�}�?vo�^{`-2G�,n�եkc��#��� ���(8�OJX.Ǖ�zH ��֥A&�2gS��,��me����ݓ4����g����h"G���D���C��`���Fq��H㨋I7��Ȳ�ݙ#xbean�A=^�#?�3�!�X�c�FӋ<�rL��n�$���t�|��h�_��N�,җ�^��
�b���{�p2sQ�韉���� %NY'�<SXv��OG/���>�X��Zt��5XQ7��2��//�ی�R4��7�.���E�x� ��-+o`8����B�^���Q�<������wOeNȞl�c,���4K� '�6��k�Ӊ"��5��x��&�556)�.�;]��fK�OФG������y7 �_��iQǽ��%�w�ذ���E� B��É��=��VO�π���4��t/�Ӕ����HO�'k�O���d����J�ޒ♫&}�='A�H|�"Cj����PИ=!�����&�֨u."�-��v��1�M��?S'9�{R�U�ag.%=��32֢��7�=/��ų�gVX)zϪM�A~$+�-uR��NmC�����V<#8�"h"�Ux�r���wF�ǈC�{�H�"�i������Xg�uZ�I?��l$'QY��^:/�x���+p�"���5'�W@"ޖ��M�(��-T�eòU������$��s��2lO��7�`l."��L)&F��{
�P�;�n���@m1'�χ����Ld+DI5��¯��3fG���c��1���.��ޡjM�Ж�.�:Yhm�-��3;��RG"8���M߇�{L�콲BV{�LtX-d֖��ڈ�L\K ��I�f��C��;Y��6����t#0�b�L�/Yω��?	^#�	iD悐��gJ�EW�p�M�D"�[�����d�C���\H�wۃW��ON��RG) H/�\��|2*�lj�x���/E�X*�h���#�j�ېL֠��9H��
��V�a�?� �Ft��.c�˥nejiҹ\~k!��#������ ���hy���^�3N�a���Eώd��Yc��8�c����/c�ֿ�,��ļ��3��4��SIJ��� �z����,����>9C��2@ޠ�I��u��S�� �|&ı�h�g�"$Kpќ�
�:V�����-�,fS��â�$�p�'�`�ehA0�8�1��N�����ߞssXc+�_����q�?%�'
:�)�-P�Rm"�|+8�(Τ���h`����\TwTY�=��E�}]�,Tz�k��EȞ����0����q٥��j����FXo?)����o�Eu�+�V�4%�rr�m}��y���¢I����������Fyyq�Q�g�P$f���ʓ>9j��E�s�k��K�K�CL�e^�<Q�����Ow<:W�v�lg����y�0��JI�@'U����WEk��Bf���/2)µ:����]kn����\t�W5�w>(���\��N�	e~����c�9(��1"�=�7hX$&9T@�Y*��� K
��2�{���gv1
��vgF�[8}�ݹ�K�ƙ$#`�b`]�Igm�dj
���J���x���(��A.��@�ɥ��(����w_Zp�u��~MuǝF�8�w`���] �1�c���Ĺ|R��q'��`)�F
��!/Len����H��	f��CD	��f��U����$�t�bМ�ݹ&���!�k�[3�����lbG�����ya'�.�c�Ҕ����H㔼������T��Vz�*�v��ϥ��0�Y�1�K�B�A�X���
ac i���Vn�(r�,���D<8[�xEd1�E��wPa���BA&��u�n4l?��;��\x�{�t�W�I/Ĵ*k �i�p���&ٱUz��� Gj��|�pF�L4|��p��w1GcT�a$w�l	b4�p�P\��]ߠ.��E�/�
�YP�7�B�;����$.��A��C�_[�Ig���H��q�A��pϯ-�༅Țf��A �4}k�>��Bӳu��$XV�Xã��'��G�SO+Ѫ��T�����K�;0��Jk��~�G����vͲ���*\Yl���T�:���m�_�a�r((�������?o#[Qr�z_��b�(w�Vԟ� �����KP�%�����b#��݃\y�$���(� j�{N*8�v+4	$ئp��;��5A�\�3��%�"���֩�X9��m�y��y�I_�  �� yjQ?�V��g�҆��cCO2
�.�_9ї�B�ˣ'r�xď�P��{�e{�`^��K��h�*%�k�j���.l��b@�C_yR_>�`�k�{�qI�cv�����>���p篴�a���ғHV$77�m-�%�m^��'��Qs1�E�S~�2i��B�؎����y���F@Z�5r��F�E��������Bɑ\������B��2/�;��;w�g8o��~�B�٦Gà�O�V/Y�y�0U��v��}�^<�y��5�pz4�[�H}tc��W��R�N�q�v�H�n|�L\s>ɓ�� �(��x���{f�mp;}t�q쿸K��Eͣ&�TC�?\4��+���Q6�����dqhoo:W^&R�:�?�T2���XA��@�3�v�����aB���^,_��8�+��_�9����Qup�i@q�\�.�+�J��̚
�y/�!�|W�r�V��Cƿ�P����nL������7�\K?���C�ʏ��v�[�r�5�|��}f�T��g�Ec�?�ys�c��=�㔋�AO�h���I�:��b��(�!��LY���5�:Sm ?-P�I<n�3��������rcCƛ^zF�S�^`1,O��Jr\����:���*��*��� ��\�tz�,�=�2�6h�ܐ���;�|������-E�n��:�W�]8���P����+�4�3����\M*�n�.���.���Z|�@i��Zc�o��Y����$M���UĠͭi��is;��c+�Ҳ�����,$7:�[x�����3Xa��D
iD����q���?�V��X�� �e�<70�g!r��������.5;x�Rx���}gԚ�DG�L�� ��%�yv�ǁ&?W�cy�  �#���/.��DdRD�%_�
2<�+�8��tG�X%}Y��T�V�i��m��}ǥ�iL�-�!7���??O���Y}k�~	�q5tQ&�)h/�4��g�n���A�p�k�KE讑[�`\l�A7r�
a���	����b%|��n}�M��e��.(?�>�&Z���SD�����+aLuR�2����W~c�o3RMYkzm''4�E��N�>y�=G/�e�+p��æ�@B� X�HƷw��:ax:�^QV*_�0����� �a���\Ar'5Ǐ0�h�D"Z��e�C�߸R��E����p�l�i�\U����o}����Ad�xw���ZE)$��,;�Ӵ=T  ����}�! �U��g�(:ڇ���lә���S�"�� {���A5ַV�uz�޷m~�� �	p�c2���~���S/�̾��:bQo���Q�R��š��00qze��GS5{�DH��GI�_4�]��fW7ǚl�	1��%.!��p��Ƹ�C���f������/䚈�X�Q{e�A-vZ��Y'�c@�ȶ<=;��L+�j��>[��)�I}_0�ԍ��!� ���Z��u��R����GSa��L�d���2����#�$��J��0��%�;�n��[�k'�����Ф��Q&;��M���Y��8�s�I�]@T�X�G���6�@}Q�9WI)��;�:ċ�dژ���~��(G�P<�BZD�G^)��k������&/���mɯ���B����ֺ�#Kw�t�?����@^���1Q�Eo�Ɣ���=�U?%���7������95��Ls�@�.����+S��9��7�� +}��t����r|�"�1�<9���T�����H*���9<���(t�wו��逢S��n͟��+V暨r�Ă�c�Ai~�7$2��\�iSs\�wX�W>N)��C ���[��r@ypa��B!$R�!�*E1S�E��A�D����Ff��ݐ�����ݚ�J�t�<��O��%�����Oʼ����JB���W�^&t��po5�u�c���ʂ���`�����O5�%�Oʴl�!z�$9il���nݣ׷�,kW0��S����L���L�1��6f��뒏I=�c�We�b�fA�a���x[�h��1�3r��k�
8;|�����TB{2� b�!`�煓u]Vc�T���-���m�!
�9��t�W��ᶣ� ���g3�)�:�v���&<jC;7�N��5~��q��� �6��'����=,9�Z��6/ �,��xa#U#BO���5�Ԋ�S#O������{E8�Ly��l>�Nf#��jE���8����>�(c*C�����_߉$�HWx��J�`?�^�o�EN(�q�U��Վ"�p�vt���?N�������sN�X/M�h��6��g���[[E��L)䀶��bkR4.Vr�!+<�m��.�P|R\�չ�̬�U�)�RFJ�[�]�gi����O�#��;�ݫ����#�ʘZ����k�/��\��{�����H�2M$Y�L��B��/���8d�>�.�����ٿ'���{cO��<�M������q
"L���t����[�FZ��fg�t0���(s�EJ`�3���{�@k� i��#g��\o���S�R�����������4Sqhr[�A��1[8�ٟ��2W|!D����o�8@<hٕ�m�r�)V@��v��Uw���5���zC	M�E���q���8{�~���b�
���`��$�����}E7㫑�EB|I��9���@^N�*�T�{���g� ��N������u6?W׳֗K������ЪE��o�a5\��٤���ٗ<(�Y<��{����.��j�z�E�t�<��vI��'�����Ce)��[l���SJ�?��z����8.o�J�KhV�1>UY���@ΉT��p�c���A�����c��)�R(%�D������n���:NL~��ҽ�}�:x�+otyz	%G;.5	�{�f!O
�Z+��KG-�䂲��^~H�,� Z��w�J�D�&ӣ/Nɭ�I�X}޼�97���{���8�᭽i�7}��o�"���i��������2��̻N:1����dQ��s��_��&���׽wa�C
�+� �K��e계A4#ŭlP&��l<!�~� �?.�Z;��r�z���|/"��\��V)<&ϥ��x�_ѻ��W�wȱ�Q�"Jl@���1���	o�l%v[p4s���@��i�����O��8r�	��{�}��'�>��`��@\��d��1m��:����$p��Uc�R �;jCC5O�,b�=1����/�1�8�iXN�@�X���A^v���X�r��.1�ǒ�Ii���ƧNG��dѷ�L���h���,�à��t�ag��.q�j�?�EQ�)��g\T=��r%F̱a8��_����~Y6mAm:��x�Q�o�8�T�7�C݋$2j=�Q��\<���v��d�'�y�A�1�-ڐ����/��AV��[�M�8]e����m�Ӟ!���-ؒh�x�J.Z���w ����� ���W��a^5g���T�6r������-�^I�n�uD.qc� �_t@��� #�<>����m�Dr��PV`�:v4���pK��_U�fTw�L
��r�%�}^��Gv��-��o)P��
d]Y�sX6w �Y�F�9i-c�����L%R��J�Q�E��YJoh��Чd7�S����#W[V���L$A*Ǵ�R ��G�`sX��w8`dck��9�4�7CB~�h����@�KC�[�t]��"f�챓
�A�"Ч���tOvo���`�i{�)NG�HL�.Z� wB������䲗�P�Q4���|Ml3a��� ���^���S�|6�82��>��<)�f��]�tک�k���c���!�
-�j�QH|c�MpƚCU��3�x��&�i��}�7 %.�w�:|��ɚ6�Oo�;Z���㭺׼��}@���Рh���P9�HK�M��ɄYW���5)��J8�o�$���}���+�F��w�\�lG+���������;�49o�����
?R0O;���B���ؑd٦�2VY~���'t����T-l2-(�\:\���{}�b=�� ��N	�!���c���Lz�p���<�cxw(�>�8���i���6 ^^y0cjG�zd�ÿ�b2��[�B�N�wF`��qb�΀`�ڱ��2�E*��EP9��o��gz.{:Sb^���elT����φ,���mUB#<� �O\�G8��Gp0)_H3�񊢙[�Rav���kP�0;�^����Ϟտ�I��/a�ì`�{�j9AZօ(�\עϽ�� 	�ý 5�Y%T���e��`FV|���ZK,�*z@�(y�(^���ƾ�G���{E��d wŤ s�6[�X�1F��Ѧ����O��xZk�k!��Eh1�kE�t��S,�����[�{�0l��Ef8R��l.��2o�bbu�g#���x��Γ��=)��xD͞��R仚=�<@�A�U QU�d;�V�Q��]2L�"�KCo�w|���Ǆq D�B��ᢋ)�!"�L�����82+#?���
�����ķ�@�8�#Y��m�O������Wb�Nrj8���� A�Q�X�Ա��3!	|�^X�]M������D��>φ�ܭ�2�S�����G�j+���C���'�^��8V"��E�Kr�cfW���FO8��/M=&\ٜs>��lY�1������`]��ds2C�_]�U|�/��>F�[�wzyA�J3�h{8Y�g�����#�H��%�`��$wP����8��"��Pe�z����7�RE<X!�pG0l�-6lSF�v�5�UZNh���������*+L.��P�f9���'��!j�n���SG-��+�Y88�dv���"x��*�Fڎ"̼�T����3M;��:
��+c�aO�5��l��nUհ7��q�Q(16��?@'���?,���1U.l�B���D��ag��B{�/�=�
�fs�N|Ze�(,��(�����ڧ/�2���b�]�Ȱ2emp&����O��5�ݒ���4��ӿ3	�;TnM�7��.��˗�T�5����&nI��n�4��9�t�0�I�lN�i�����>��3٥�)��:.��S�k��T�~�VO�1Kׅ����ͦrW��f�w�g-�f� �Ps�or�����5H�>�>�Cl��ׄ�I�'�,�M�B�g&%�9��d�D����Y�� �(!��|7=�V���ޕ)�xo�M��vg�, �~���?�'\.$G;���.�1��lNZ�����K�ر���
��^��gn#�)Y��#m�}��F�-x�G�.�u�b����ˆW	p�!ԯ���A����\j8�r|X�p�`��|���87_��(9�/1nHl��"��V�めW.�`JGq#j�PR*2�I�L���FHѱQ�fm��^��ܠ�d3�.\!7����3�ڂ�I��΢��^n�zS��B�ּ��</�I���$[S�T����Q8c�B�0�ZW�7��R3ؖ4��[v�JG�ä�H[aPn|%��ë1(�,�l�@�p���e$[�~x"�������[�i�z�((;��gp����pb�d�)��䅢p��j��ߎ��筇���0#3.��t�2���ek����{W{�l䲻ă��k0Rx�T���A@�s �\DH`��%�(�:˶`�?�ҡ *.�GyxE�r�C��K��������v߸e7�  �I��!����MzͿ�sDp�B�u{x���[2b�S���/��ZQ�$�س=p��e�-��m����7�~YC�|�E>~Tf8H��k�d�|�J��F 8��}��`�������	I��t$l?�ݽֺ7	���ee���ϛ3�]+����D��O����f�OGv?�Sp��P��Hu�K��3���yc\$�eOB�Ii`��uF(�k���'�k<��n����e�H3�)�,5*�ҫ��<P/Wp>{���W���O\�G:/�q�O0�EW#�i}��ܱ��b��8���,����S8�Ю z��%�$�/��{]:�I�C���j�فn'��#ܪ|#�m2��ӳH����0�
��g��zcT�O�@S�"�o���]JiT�\�t1�]���e*�"qu�{5s�+P����'_V�j�\I�k��F�S�(9��ZѷԊK�8޵�V�C��("�y���t�d�΄Z���(��M����C��n3��{��Mp�`���y8�b#�X>�g
%~׃3.9ݳNiR���I��g��Pj�b�_��[���<�� ���h�,G�)oE+���[<P+'�(J�Մ&���2@�.�uMvw���a�%N�f��c,a���S8̸��,�g�N��]�
[�q�R���gK���̜#��	o�_ s�|���һZ��������=)�V������Pd=�~�JE�=��TJ�C���S$E���HE���Ngdji����6~>�~\�*�JS�R��Z����r��2.���w���n[��\*����pJ����	��v<'�n���������J��C
4jx2n���NJ�'T�=q��[�0�_�FL��I�7U�lϬp���F�lu����W�u�WR�E�������O�(��0��[s��#n�F!��ا|�p�%J��į��
��	��6���A���C�K��P(���ї+%d3U��z�J?FΌ�xm �,(�r]v]���衕�גZ�þ,-~F���cD�ꏴ�S]Œ+y�kR�^cg'8�[���b�kdUB�m���}�f�]�����$Jx�ƪ�]t�M�N��~�~�"���r��\̂�i�5CXE��OG���H(�	f[%�O�-��Q�0T���&�����0�nRX��������p��^�P�j(�-!��f�b�OO�^N�'�K�����ŭ���)�=�c~)�=��[��2�������s�G��7
Je}�8�q����ی�;����{��~[�T�P�7k��͵�Z\~�r�8:��[4�oͮ<:=�Zcy9;5g���d1��iP����􄟃}���x�[���\a��ީ�q�:�JP<sp��, ;�Q]v��]`�2�>:V�~�o(w:�
�A���bev���4uP̢�o�QbW'=�uG�Qs.3V܅��q����"U��$�t�RC���	9]�=�g�:�^H���E@�KE�7p��$��>����Su~��L����'&��,�} ��(�z��g�\��6<+���:0mҏr8g�ɠ��I}i�!�@9�u�#���Ҧ�맬Tp��}	�C��������v�*��2՟5�����$R���_��Ar(�ج�������S��6�=��!�����e�Ate8������p�|�f�2��3`�8��n>ޒ�D��9`_��;�Q���Uq짿9����1T#-h������
��K�"�����N/ e�E�=YpF�$7�/?b(���x*J��&dla9F�Ö__��	��^G]�a���<� ��.�3<K'��Y@�{�b�ĜOϰ��*�y�5����ʐOv�6Z��\*��-���2D���Y�<�.vf��x���7��[iX�/oPu���y���᜛tI�w+̋�d��$����w�q�>�BgZ�:�[e�y�\Xt�+#]�wɦă��_��~�TvAo���� �j4Q������Q�����P���cQg'F�wr?�4�_���I�����g��1�bmXv(�n|y*Q-�A+�����j<�t�<�Z��wg��G��ژP�yG?t��&��Px���s[G�x� �V�um��ozł�)ڳt���G �D���D�V>�*M�!��Ώ�����>������4��ڝ�$0:yo6�� D�@~z����&��"Ԟ��{��!���i�N�5K2�Ү2�!A�-QtG؍{<�+�_R�珉@~�U�ǶA��/�g��P�-�ST#�wL���?6��R"X�S��R�K��b3't-�<�eC �k.�Tgi2��u-)%�Q���#�M2���H��kCѲ�S��.'qQ�0�j������ ���u��L�_��S�$�]��Z��oߤ	O�ӊ��*u�����fo�ٶ������	�s撱nK����Y���-����ᯛ���E��&�q�f��~1��`g�Mx_�=ag����2�x�?fx �B��&�A|UyL�^�Fئse$Q����T����j7)��u�ײת��[5ܟnB�}7y|u�w�G�f�n˞rXHO�΀�8H*�����we���Õ�/��1��$J�߯2}H�8��C�jSʎ�l�ݱ��I<��X%r��⹡��r��E��������)Y���l�WV��h��L�LPbd�k�SnS4=�nU_\�����h�Q��?��"+�1é-������[=P�U��Vr;�ّ��=b�N.��E�6���aɠ0�Rȇ>�g$�TKS�k��ظ��`B�*@�}#ĥw�]R%/�땕0�c�.�A	Z�Ff����-�Ͱs
Ъ�[ZOeU;67U	���d�v��A���y���e��ݱ�+3�v��1���2��2%B��9oW7���>�9���L֢8�VX'������l��lcE��ʪL�Z��Oy�j���G�RLY��UL�&����*I
��?������ߚ��UO� c�hxU�s�4��8�H��V_ji>�d[�%�CN�M2�d��P6���8z!�x|%d=�ۗW�G��-n��8V>�y_�l/�Vtu�Lh7�l1��y-)&d4�/l����a�F�&l���H>^�s�xJ�ѺL@��PϹ>:��Q�Kū��}�D.`�-�H��.����[�����G�q��!��`�:��e+��ǁ�����MB�/J���
�L�A� ���k$�3'��t3,�[�8[޻M�Z~�(���,	��l9ⴤuex�P���` �^�[E�ؔ���=�URM|&�X�:����jۻɹ��!,OU��� ��Кbbq�0��	$�]h��<�v&v��(	*��ʽ#�Z�h��U���"�x�ܲ�˾O�0yl}�T?�ů%��S
)�tu�u8�+Sހ����"�љI��|QŔʹ�y�C~r(#o"E�	���&WF9Y���}�V�#�B'��.m}w�)�]L��l}/�Me
�9m��VF�s��0$�,p�ϧ�ne���S���1N���?8 x�?�W�x2n��2\�8�c�e;O���,��~�6�<����io�j�M�޾�G�	B�ۜ`�ܶ^C�,�yy�
bd�s��r�$3������׀�qѣ�(ΰ��� ���:��5Γ��	���-rc��U��P~H�T�سp&D���`N���͇oI؇>M�WL��*O9���<�������\[vF���(.��U-IB�S�L�t��e;��r
�	�<�:?u٣F\��q�HY4��6~+!�hjO�c�0�D	j]-���B�����V�_���&h�8�=�1�Ԟ��s"�cl(�=�{���� /u!7�Q���_�t�[^
5N����yD�]#�����Af�̓&�F,g�����f&�	}�-�qy�%�3��?�`x�*-���C�g���#� ��3�z��W�d����5}�x�ݍ�5�����]R�f ���!mYW _F�ns�]Dt�|��{��(}<c����ۿ;�U�L��g��m'8+n�j��y*#Zh�"W���S�U������ӎ7�(��p@{AA��T.w��C�SC�� �ϐ�Ȩ|�s�ہy�R�8�r�Oj��6�)�wgt4��QS����y�2�A_�j��]�LZtp��Ck�5�ṫ�k���`��mFf��������6��E�ē�ړߤϣ��@��:��揎SB�zZ�`]C�5	n�B�{�#�M��Ňʹ�V��Ww8$RV+D��Bk�,�	��30����9zڳ(���\ysWJi�ux[V[���p�����3�t�bQo2sq�zA^s��К���qcsE��' �<ga�u^��y�k	�����G΄�]����ʽ�+��F��P�C��Ճ7Rn;�FCVf1�s�fZᡘ8�丞�Pn6�+��E/R,3���l��`��<�2�!'�:l,5�u�0~�68��X�ajJ]����#��n�}�|j�C�#�ټz�$&.���G���)�� B�3����'&��e.Az��R0�c> h�C����1�_1�3km>���P�ɇT�^�:�i�X�C���-�!�0�8Z���&�D� ��$��=.]�b�r�'���:�uޭ��|8B(�$n��Y*⩊Z���G����ч�އ#pY���˕�0BS��fV#2Ot�{(ܐwmP*��U�e0��o-">�;h����gv����\3`ޡ�(f��$uѱ�?Z���"�Ǚ)�8��!߾	L�M�H�z\��v>j�됌�Q���R^��Vv�G��j@&�Y�A�,�ڭ����-i��jX���J��Z���G�<G��Ӟ}��[oؑ��G�׮�YN�����q�<����gd�~�,��)�J��7�jM�~�����56��/���9��τ��K%X#��x{Xe09�A?��Z���4r��Ɏfe
���)�)�@K�o~_��$�7j���#��"�F����R"�*���\k��*}R�5�b�O�k��Fѕ���;Q����}{R���H(�����{��=W�t�5ݖ�t��	O���H@�-�ȯq���n���-C_u� [Ul��c0���C~nF`_��g�����Ԣ���]G�҅��.wxV��T6XaG5Ԫ���CK��clR�a
���Ĝb�Er��	�o�mu�R�e=\�n�%@�)����,4��3=��>��jV��p��/������M�ma�������o���س�bS�\���90F�S��cK���6����m������9l����F	��Vj�q��(B(�A�_u��:hWN2�$�A��g���4UT�N��q�P&HWh��J��o��"��_�9�N�l�Mz�(���h�T΅�V�C�C}5K��F�í��Ӝ��I�=���_5���c�a�m{��J�YT&�w�S�����z�Tj�,B�q����I������Ib_�Ҡ�7mB�ڔ�TR�-r�!���jL��Wֻ����Q�<ԿG,�궾 �On1��uW�%kڀ�i�� �t���V���\�kC����<�-�$����pн����%LixeF�YD��4ЏL+��<�g΃���c��x��ȕ�S�������:�K��n���WϷ��p�df[6�����7���Ob5��}jy�T;�׍Dw��ϙ#��w��pn�&��4+�Cތ�}�0"���P��Jo��-d ���w"�/�x|8+�쯨.q��ƪ�Ba������+a��qX���b���Ll~FάL�e�^+p�#�o4W���KN�����7��"�.���	d��)I���Z}!XF(�^��S�s�HB�� ߟ�q�P��d�f;�v�_{;|�xT�T�,�i��e^ZV��`��o6�3r��oF�a��e0�����n��6g&j���Z��9�L��]B���Y�\��:;���Y�q�o@�'�mZ�js�f�AGH$�ڙL@3+�x�-�_'r���E�ۄ�9tT�*Fv�%�29s��Z�����+�ׄ��`�6�E���͙1p}N�EE�50��qI�r}`݌���LBwu���{�����֎��Mӹ}�Dh�����x9��L\;eq��P�(�T,"�Z~���5{��?�\U��7��y<I�����,��U��H����g���:�k˦����@%����2B��+\��崪p���CE��0Z者Z8'lk)&�͍9��?nM��֪x�&��?�1���?�x�!N����=n�%�EB��ԕ(=�8W��Z9$,���z[
YQ9B�[wyL	�cb�����E��N��Q9�sE����#��=�0J�["�)��Z��O�2?W5r:��79�Ɨ*�4���bp�x�c#�z4��$c��J�kh8\�$�����x� # k=�Z3Pw,-���t<k���/��g�ok��Oۜ�>�KD�������� AДR+��Q2�ϖz�{���g�_ڝ���J�`M���r��q��m{��d p�+����XhS���	�'�I��	JD�r���d��ȹ�`���ڞFo�+�k�2'�������UV�TWch2F� u��4�$!$����?�!�K�-�Oe�_6[2�[��yoB$	\��bOh�K���̺�N�gdT�
fE\)r���OdM���ժ/!$�+l��7���}m:��Â��BR	4i����`�YT�p*邞�g�A\ř_��h���J�2�]1��{^���_!�E�k��Q$\�i�(. I��e�3(y�|Eɞ\¢��
(%a
~��Qj����˕���
�zl�*��3뜣i�"���D��6�?�C���c7�"܍(mo������z���m=�=d2��|o�P�
=��n�LsQ����,1�$L�mznV0ݷg�j��w��)����8Mk���\0��;)�j�tt�x�bP���2��k���o�v�����$��O�/�Q.��� ��G��okd�Ƞ�&�=).���n�I�>j�<�ݬ�0�6��Iz�HJ����݆S�C�NY����S�V+����^����A�C���wڛ��뙗�����,�|C�)٥��O��m�Nrn�W;}�Xh����{Ní3x���_�3��aE��ؾ�i�n��(�t*� �����ۦ��>�9��ߩ��R��j6�DX�@U�T*Z�_D"�JV�Tz���\b��6�t
�Ih<VI���4���ARn�{����*2�[���w�ƂA�QX����챫���Vr�8׉�ЈD`�UU��i>O��8\��IU����~Fh��{[�%ev�'e^:?
��Jy�Nv�v�4m�pY v(Ţ��<wye�h��Q'Dt��x���d�F��" �}��‵�ܥe����_`۲�صl��gN[GLG<��:�����0GҲZ�d�x=|-p�[ʻyr̋s�����w}�w������~����B�o��V�U�mg����Lw� �9���`�ՍpH�����ɇ�*�M��`���O�*�4�n�Z�ݹd�X��W9�i2���^$��g'v[�_��6��2h7=%�����).���;���g����c�C!��q��#b1�����6'(`�=�-�!�g�V�����<#���@�紐Y_����y���<�����3�4c���*:H�q�3Ur%����ޱ���i�}���bY���m�X��=�o��lY�;<���*�5.�\]6�U�`}ĥ�� ����WY&�ǂL��-4j�^x�d��N�G�k��s�G�c�*l����?��Ց
�^����'��fW�$ �*$H"� .} �pFW��ӈ�w͓Y�tkB4����Nvf�v� ����[᪶?va$�m�]_֛B	��Ӛ�[��w���2T�~6`���F���J;_��c��}���-c���t��H�)*Hb?���t��s��~�^<h?�e��̫�[T�E�_|@-��~�B�����I�rh���:#W�@'���x,�b5 �Gٕ���.	]���O�FY��SbG.��/����?^2�M&����!��z"J�M?�L=���h�ܓ�m�jn؃�k�j��5ONO�(Fx����A}��UsZK�77���c���I�ɚ�{O��?b�m�Fr��g�ƑG%���#6�vz2n|:&LGF;t?9�����̙/x��f�zC�ߵ� 4��ɟp��X�~������������-���Q��.&�����
��WT���D��$U��x|ܸ�Ԃ	����3�)���� �����k����2�(�p+�k"�̹D�MU'h��͒��=�3���f[t���6R$�xr�%U[��G��Y�u��צI��}��	2��d�Q�I����i~��\3��'��]$�(\��|�>	YM��"�P��1�au����d��h#��+���� j�o����A"���+F-�@��b����<Cp&/]t�l��Z ��X)i�i2w�<���q�k	
(�S�)�M��¸'�v�~�6�]蜾�2����\�N��"��@B�f��y3 ͐P���rA;���f��4��R7�ڃ�e���a����l�ZaО�S��(�\�E�],C�[���uR0�N�e�ST;��h�!�o��p������}�F�Efp}��b���;|z�8*�.fg��=֜��嚷�Cu��k�Qa��*���@�*!N�	-v	xG��$#�{��v�4�h���qs��[n0���Ё<e4����_<���2,Zc1Shck_^�K�5�<L�8����^��6�M�؏yω�$�xky֥�Yd���F��n�4�6�QH��K����;�N�V��n�Go�v+�G~������:��ɯm����o���e(�#����gP��ķ�@EPA� 3Lw�ݎ/)]be��p�5B���"6���+B|>o����g���d���LjJ����rC`̒�?�@D0��"p�WX��&�7�au��,ѵuk��Z��@T}�Ң��CT#� &��&�?Ś��L~��.�O�r}�J�XԿ��6�6Hk��)��,�]+�F��ҡl;�gMN���>�B��?q.d_e�i�7]���ז�1@	�aԊ��0*pg�rQ����*uW��<�����,�?���o�h�������n[	 *���E��5��:���3F"Z��[��{�3���)QҰ���-6y����a���N���J�jd@h_��)/ ��ч����h��j�6,DS{���1Ωg��j�t^z�w2>?�+�3镉���T<y���j���qN�<�\�B����h�r2�����z���x�6;���b��="�GM1L�i@���8G%�E.���X�N1�a�Q&*l@}�P���KP�w����u�a��ˆ�-1�z��/@�v�b6-uvGx��O�ǘ|�U������Nk��<�ڕg+�tT�
�;���9\�/:���p]�98�:���U��-�Ҁ~k��ׂ�̅����T(����U���$ȳ��h6����4˼����,�$!Ғ�H(}����`�q(T��K�H��Av�y2V�;�gh��O:	�.�gC�e�
7�����wuڪ���5�n8�0���"�VŉԦ]�D����|)�Z��F\�+��bo�C�I�.�����	�'�6"]Y�<nx$�JR5����֩0S�-}�|�9��	H�<�J��Ѡ��B�!)�֚!���8���ڄa�-���SfR�4��Qi�$q.�>���%V!�����I	��WW�D�� ��y�r��R���9�Q�����'���Rw����]PGz=�m�.s6�,D�q�����9��4����lWs��ю����o��Z��v}�z2(� ��/�%c),7��δg�j,��%��!�\��PᢞX8��*��
#K�=�nB�b��1e" �dKI�h9����J��<�r�} �rY��^�\ߍ�1H�u�xJo?���g_��]���L��8ad�����99�$�=XS�*����c��e���D��UA\���L*�08k�(��[�c�d "�d�F�{a����G\�ܑU�K'P��������Z4��YX9��a����߾Q���3*��7�Lj��y2ۃG���n����,�1��1Yc�v��Q�@�P���P�(�������&��ަ\"1A2S�	���F}/ �O��r�ʫ�:����Ί|�Ž	H��<fP��O۹nj�r��0��I�U��0���[�ط-�;Ws��}��F�0z�N_�ݮ�[��yO�&�ڂ�׈M�� ('|�)��_#���{k�YC��8�Di&y��S�Ʋxu3���?�"��[9�;\�J�?(��Ц��l�0?D�J)��<�������<�5/o/�}�jm[+��$~�Z3Sr;�Pu��Y�����@��{5U�n���}	�$g
�Δ��GW��'6�T��SS�d�9�3��\�4O���1O݄�3��b.Z"�}�6�:����Wӿ��; QX��	�d���<�ZM��tI��Ռމc �:�Ī$)ߘ���|�mj��[�
�aa�MD�U�g���R�Ӝ8�^C|�>[)��\֗�r��<{�#_�� ���W��|.�M�������eoG�1U�����:-?<�	l�����*�A�K+(�/����63�lڬ?���h1����>�7��0+g����Ѷ~e�j C��\�ʦ�N�AUag4y�P�5Ɏ���(z`t��2}��N 3�XYhۋ �u��ㅳN�
�ڰ8 .i��wd�I<P2��uG���� �۱�.	�8��6d�9s��b������6G#k6����2�5��ࢦ�'�ɯ�T�3T�ҋ�M�^�DEnJ����n��H;�F�5�c�� mH�j�̧i��w�tYb��σ`lugۉ�Ma�C�m* ��JĪ<�a٣�k�>�X�{1ׇbƪg�J�!��3Q�:w��G����a�aOφ��h��.�B-m΍o���v<�r`�����Hi$c���i	I9���<�f��|G���$H��
g#�N�E&��C8PX�q$�x:��0_1�d�Mx���������� G[.s�7���-�Ce�[����_��R��A��%)���B3��՛���>�%��Xw*�SrG����%�6�|G���N��!��Q����(DΏ�Ck�m��XB��SR��D]I���'�J�F�,!'��S�D�b��U��Q�x����EI&��(�~ì�3W �]�Ÿ�pO
���<�1�Zj-������SQE���q��Dy)&޾�9QK|�Wx�H�*]B��A�a\C�f�i0�ޡ$%Ym�u���e*� FF,[�����������ʍHR-��;+"qh�ko��/tє�n����_�x�������Mew]#�2��Mª������,q,��t�s�ތ��"����l..�V$M�j�%L��C܍iӆ���#a#���-���Q��W�T��v�;�KF�������8���'mn�D��'��-5*Hڂ�y���q��n�oWe�)~��$�n��+t���/�a�p�wy�$ϰZ�U�,S��(��E����ŷ��4�sp`Ph������"��M��?�J�I�f�&m3�1��|k���nG:��:ST��V��?�j��J7Ӻ��j���@��LU�˚ �c�:�s��邀�No�7���i�v�q�jl[)�)�#�"3
�r#`|O>T�ɪGo}KG�����0�=sf����ׂ�B7��
�(G���#�i�,���}�e�f|�/[����\FN�<E��༔_�l�D����Hd�_{�k�3���ĖQԘ�~Smb���ʟ:����u��L\ո_*�H��F�s��FK�)��ɫ���1nM@w�$j�K).
9F�����o�Q6y���lc@6�j�~����y�1�ss���3r�G��rPV�p��s�����b��Ċ�%��m��/	�b>��2�� W��}oV�0+�p�|C�B��}���Q��g�g��� !��.|E��w���Ҭ���������T$�z�u��J=Iw��!	��s��`G���C��RV�C��FJ����U+�p-K0��� ���k��������-����\�W�)j�Y�B���ɲ��l'�y���YBV�r#@�	P�f�bΠ^k_�ڦ�����T���1tp���t�|������)RK��x�x����j=�%Ë
u���`cG-W�͌��0���gG8"Ța}n�.�(�g��_�歯%�a�s_Il|F��� �����tI��:��Ш�%a퐤*����S'���a�V��8_5�࣡s�YS����_AG�=��%|`^����	�Q�W�$�=�,��i:H�Y��F}���GP4�1���*5�hkn�'6���蝷���v�g�O���X\Gt�q�ݲ8,"��y2~)%JI[{I��|�`�|t5߷S�toP0�|?��c^s�=�Έ$�gl��r:����$ϣ���ƌW��	��S9�<�h
�����eGM0Mqmz�6��#���O@4��W���yy�#�G)x>��M������Q�E�a�:q��o=$m�\1zL��D5e���>����!�������~�ޔc��%�K(�K��?�:d(�sg���)��Men�_�~
p��/f7�1�JQ�$O��ǌ_N�A�rE�v^Ѷ ��n�2uz�|�@#�<L��v��)s��Y5�Fdzׇ2TMT��ب��8x�3[]G��|�7��e\���^z���Ì|��|�Ԕ�$CMT� :��V�h,"�gA�x�wKf��Kr,��2���\��ė��:RelZfX��m��K%f�	p�<��r���k�T�ڻ�&����h	(�U�t��V�.|c���H�?���T>��R{+u<��)�	jE��܏���x˼(��"B"��ʡ����?��C��F�آsidA	«⟙d�G�MGS��L �{�@��N~KL�B[��̪��oǘe��^V�df��v],�v���	�C�1���<�
�s��͘A�u1����	Y�jĦ[UQ����P�ۜ��|E���hb��e9ߓ_9�+���fDm-��傘�m����J�ѥ���X�$��O�bΡ�c����� ��O@�t��"�y�?�{F��ؐ~��(�
������JS��_{J3<X��G��TT/!\��Md�������|��a㡃�}��%0٭l����8��]��DH���xB9����\�׹Ȏ%�\����M�ԇ� :ƞ|���Ҧ��+]�� ˄��x���8�c��X��9�zq�k��s� ��'@mL�z��'��T���j-��~&6��[���+5��Г8D�I��%[Nt��=/����2Q���0�/p3`n=>�|ZA�G�ޚyyh�p0j���S�}6�1��k;��HbZ�Nt >7v�������4؉w�񃢉odȎ�s/j��"��Z�ך���@X�tF��hè��Z�P��[��V��U< :�د[:��ɼ��(��pyG*晀�S���O��p��e�Q�I#X f��l���"�r�P�{�C�Q��l�zXA'�7�
��R�ͅ�b�7��)�s�3n���%a�@��ſ�{��Ea{��b�PH0�j	dU�ŭ%�kBMR�L�]�aA	q��>h؃��O��W_U���m;QnO�	��{v����	N]&���1v�UD�(�v(|E��7v�m
rm�E��(f��su����7iޏ:�f����Հ��K5s}K[p��'a�?Z��6U���S��J]Ս��i�BK@�����3e`(k��r���&�W�N�����9
�p�e�"c�b�נ�f�s�t�77��:b�Wa���aJ�����Smbp�&֮�`{ġ|��#w����a@8� 8 *�����;�̓7&r�|~j����b��:Gɤ�l�4E�(��U�|pD�x��I2�ζ�j,1�G�A���t�
��y��`��\�����}y漟[��&N%|k�}F��}�v�d�h^��un������3 5���$t��΀K!_��Y��� "*�~j?zd��I�(����:��gM��?ێ^	�#ʵ�e���np�).]*8Ag��ͦX
?k#��w�z�z�gǩ��2i-Z�R�k%m�=�X[�1��#��T�����B��Q��]�����P�a����R���q;��a3�3�r��P��p{�_�g�� �k�~3`[��!�d[�T6n��f�6��r�ZM8uŜE�X/Y�<c�N�1��Np�V�A��s�2���v�kX.���c�P��7Z��!���Q�>�V\�h)4D���3o����i6�f���j��L�^����mȪ��?�_���WƗUi�`o%�ƚ���{��{e�Jy��C�X%~�I�M���g��GA,���OxM��%,���QT<�#n4�J|h�72!O]��Mxt"����!ZȔ؃����K�K�_c]1�F%�+�@�������v�`�f�ppV���l���2�c�� �\��@X,��w8]��%׋$��� \K"gv��q,��N�r����Aտ�kb�.u��:���߉��ӭB>̂��T�L,矍
���nO�6�m'���N���_QmK��fӘb������z���.���t��Tg��� �{MJ�����Ҳ�7�m\?������w<U��lhu��(����۵|AG�"�K�0Uai�P�u	�I;�Ta�%2�_fE���-�	k��	��I�C�s\,F���5�������<C`�Q�'k��H��I�OZh��e���3�t*=��ϸ�h/O�㶗Z)�XXy&*�>��V�qi�����(Y�|Xyl�^�Ry��<��`�w�����WN���tʹ�W������4�x��$[�8Ek���_j��8i:�m��T5Q ��+� k��p��6�f��t�^סn��%J	݊ �7U�)�{��r��>&z*V�aM�Ō�t:0�I�_D��n��"h��%��~�d���_��a�J��1Y�M����ûG�RZ�����4�QP�Ѣ��&3}�#x��_ߜ �2�z��5���l��:�e�T��M��
I��)�L�"+� ����=�+���
�T�/[�a�R��n�&�S.�B��">r�&y��Y��ZtJ���c������t�9���ǚ�ZN�����Z�zű����'1x�����q�\��������qV���nb�U�F�(�������#�"�ִGA��5᎙%�\bᶺ�7��#��z3\V�>����$�W�h�7:b�t-��~��Of�-VS�S���Sh	%�[R���+c�����.:t�5{-F%��%T�;��׃�e�K�I3��1&C.+~˶���F2�-Io������\���89Y4P����V��l�jp�k�8 ;+r���F����&����yY 5<����l��bz�5ُ����*"� Mvf���[�)3jE�K?|��T��d�>��h<��?[a��/ǟ]�����m5����j�KU"cj0@�2�Î��l�l�D�\� 	�V�+�����ǽ(�&AWY�@v��ќ�� �)�a�J+�h�%8lw@�z�è�T���s��2l��CtB�0y
/I���������b��MZg.�٥��Q�� ������}��V�指� �H>�@�]���g�[o'�_��n�>].Ȕ��*�>9��Jx�~�֤�b�� �t�X���Y�[ET6�A��%' t����µ�%	��=:)0��HL����[���9�80��{�B�f��h��5���Ώ�{H�S�#,�
�UcN��D�){�V���":Q+4.ޚ}6=�g�d��yC��\:�˭�S�5'�}vb�΃�6���+��`ұ��v��(��g��<	���U<Δ�ɣC���Ҥ�K�A�p&:a�����BF&���6�����r��ׂ�j����>P��3r׉z�ᾗ?����Pq�o�����˗��"����XC'��̞7�ۜG�wX�e����HhQ���z�g�aNrn���NOM����y`T���@�6uL ��w���Gk��X���ڜ'q��]�ÿ$�*�?�ĚW�Հr������߹���_��Mߝá�]�%��@M�?$%���O.: a����P_�Nɫ��\�IV�43�f��MmW䞽9Z�9���S�-��Ғ	�7��A��NL�-�R���u�ir��^�MV�t��y�+�+��EU�lř��U��,:�&l�Ga+�m����X�op__D�t\�߾쁈`�Q��~Yɺp�O�O�'y����R�!
 �ؓ��W\�#�mt�S�<}$o��x���Њ���G ��
;� +￬�F|:[��F<Z�|�:�ن�W�Ϲ�=�߯�(� �o���Ն{����Vˣ�A{UW�����
�g��y�����+�hOA
 #5��о2���?�&1�__��I�F~�t����T�(<m6�o�=�~(�u}��bqi�\�7�?��G���[uh.���˄2��7��h�[��2���հf�;/�Jg��|���c�vK���xx}��߃�Q����Bg�M�=z��
V	��C�Sl��xB~A�Y&�Q��b�Ev�W������?eG-\*��;o��n��J2���"v���������&M����͗Q���F�'U*΂�&vW/��u����
�xq_�6��B:8�~3���I�q�%���X�S���9����`~D�}V��]�:�-�����̱��Y� 80�n�U��=�q:bZ6H��&%3��!�w�`�}��y�rf-��|�:�"���s4������d��]�\m����suBp�	:���KF'c~k(Z���6��2i����\L-�|����`��3XP���<km�:2��_]�Њ7��	��E�✕9���ݚ
4?�-,#}`�> �;��m �����f{G�a@l�ݍ����;�!Y����%?McF8� �A1��M��l�Ew�u��d����j�N�Re�6�Y*��j�	p�k�Ӈa��B�p("��s ���-�XvoD��K�ʧ3���_�'��F���]bt��cY�l�ӻv��{2\)o��l�z�<����å��H�hz}��:?�\�01\���m/k�7�L��纛{�<R$��γ�u�<��5E6|#
�3��X�AG	���ZP^H7�iI\Fі�g�_�Q�yR����^�g�3����)�d�0��	
G��]�k>����sJϷ^�&0$�[r��Lk/.a�p��'��{�1�&w�9 a�w���ω��Lq��|�!M�ĺ"Z���^�Q2}�aǱ|���Hry�ƈ���^ n����-�W�	(�)Rv�?�U��8���>�k���6���3�G�_��sd".u3��*����c�it�Ɇtz��S�g/�պ��Cw2��|��
�1������`^��i�����s��G�2���Ewa���u!#��<��ᰛ�}�!b���eU'��{�i�cDB�`������o���/����_���C2U�VF�3��U�76z�y�1��4�P��n�H���� ����Q�Y=Z@٨IP��A#�N$���껧��8Sܼ�(�7�^gl褏DD�p�i޻j&�LV�p�w��ܨ{Zk������Sl�t� ��\Bcd��0>L����d�pt�f�I����P�-E��k�*�q���5y� ��~F�&��ׄ��@Gp�	t�_.����J��ÿ��]E�,E�Y5�aǠ��8.�'/����y܍�>(���Xh����,��	�?v�[~�$��:<<v�Ajʌ������zqy�����6����7��~�KR YGû屭�h�APB�����"� Ke`�@PD�� `�w�a�b��İ�B�g��%d�o:���(SǮ�
��<k�m]]=*��mL�-	#(��g,��/xu���60�51,č�m��Ļ��(�TSX�
�i^@����'�Ź%����A̒��Ч|�ڷ�+����p�Yv�g\�&���^�,�w`%l�P���v�$U��Ykco�f�iq@��mA`y�E ����iuZY��{z�"�D���v����ӷlI��/Fs�����(7���p���J��ط�%-����&� �i�v~�U1��L�����4m�SqU����%^�<���>�!���
<F���b��PP�2�{^��Я=�����N~
t5�w��.2`-�����8�����S*j,����I��+U����W19*�	�[h���ݒ��l_�
E�����|3�=)ݚ*0�W�^�d*�g�v�{�����	5b+�x�+��U.P����U9������H>�e^	��t{��a�G�xz�������x%֌�Cu����-k2��W�;� ���O]���E��i\�p��&6�xY�ߨF�`�l�z�'�Wz8���)nG�UW�fM��a�Dv
������[2�$^r���F��I�<�9ሖ�ǃ٪Oc�8�٧�Q����"@ ��r��tۥ!3]BqJa�c�:W��
WWB�[lI���P[��D���m���>�L^e��ԵtT��Y���e �J�D������+� �(*xTޭ�T@���|�V|^�Z�b%/��毝ߴ8�G�&�ߵ����"Ű�6ϩCq-�)�}x�3�G�q����}�n^՗׸;B���Fm�2p֤��*h��/�K	��gL�K|{������J�l\�a�r�3���ڇMp7��Y��)����~GR�8_G�i������X=��4Ќ��ȕ������� Uo���A�nH�p
P��*�bN��.���^�߄�B+؅FI������J�@� е)/�g�p�tߩR,.d.@���-u�H��
~�3�N,���L`=M ��G@ҝ� q���8�6QAO���M�crq���oM6a�i����uQc�U81��W$�)���}!�[N���=����\����B����-�,C�{B]����n6?��/Tw&�[ا��ʖ�p~�H��|X�0'yak5��:x�ؿIe]g��l�%HK����`ҟ�#��G��]b�����%�2�L0�P*}2�& ��
�P��ݢ���@�\-&�k]�����ֆ22TG��qq�	f��hg��*y��c2���%̒��ttw�F�ƙ��α<�����Q��M���A)U���y/uR�D�;!�b4J8+ͥSr�O����'�E��p@4+�C4W�z*���)��X�V���WڗL�L� ڶ5�Ȍ��!WCg,��G��q�M�+�H��N�E�h>3�1�ڭ��3����veX�C�Ɓ�{���v\�0@.����s0�M����^��rb���pS��1|�!Xe}^���'��[=�'κ:����9��ѩE� ��=�+��<��B��(���Y���G�%�$%����<a�����.yyIS7B�I6�>
��'F"*�1�#��ɻ�Q�`nд9���G�Ln&it<<b�C�W��h�W����i�6���5��rd��x��$Q�B=�I�\H8Ƈ+u1�%|++��y�ʶ��ɻ�V	� �C���!�ꏄ�r��m��79=��*n�xd���Ok��~ݵ�{_�b�m�1�����(�v^^�M�ء�kp��c��׾��S��_�#i�KZ��r���q���+"o_��x\��@���-���qaE�<�m�$�U콽�Q�hJo�W�1�J(�����i���u*�G�t����l~�}�13�Y���a$��%?^O��'�=��a���^⑪�^[8MXp�
x�ЗUө����]���!=v �R�w �Ղ��#���j�e���h��j����(�PWZr?{�7��hfp�OH7�������*��+�j��}E��;��1v����],�O#��t~Œr%����9��9Ԟ���7}��.�b�Zƿ�(ɚ�hE��E(��RIy{�B]�R��!�V�.ß+9p��2	&�[f�b�,���-5��\���^�G���fD����_�(��3N��^2���Tl�P����N���yQV�[�?,U�����eI�Ux�H���[%�|.�➖4�[U�"}%A�#����L�!G#͜���A1�[�m���$B��TO�	��N'���΂0��?���|#Lk�ib���
a���w	g�0����6m5*)�8P�]��UĔDi��'���ۜ�* ���,>����v�#Pl'TM��f�=������_�-��?��m��5Z���rO��,��l�0�Мt�v� #�f{���0�� �#���ӗgWFN�U:"57��U�IQ#�w�6���-/í���-�0a<j5rf?��Gx`��}�W��eL�� ����ѱ�����lH����f�&�]cD�v' ��Q�+SK�na:�շֺh�O��ʴ�׽��k���+|����5㟔&wy]~9iv�)X��\�Ff�*Lx�@�wf_8:��e�}%+$?mb3t(����X>�"� �����(�SW� �K���-�� ػN��c�?		���c�r�Ы��,�Sy��i0�G&:QP>���AjO�L��z����,v*9d���$��kY��*7�u������<�~��	�e���i���>������뀸�/s!� |�5�]j�mzV�A(X�����XB�x��T�����n��:�"a�ֱ�W0�3I�e�E�����t)R-��a��Q������hpD����b�yu��cc�n�!��i��d9�VS��c5��ԹuN�4�D��,��0=(�[�o��(+MZÖ�T����ƽXJ���K��T�Q1U��Be�#�[��RE0%Y�����ȔVOH��a��U��<�F�L�^>=�
R>ǳ� �U��%��}�K����:�q����|������%ẻ�P
7����������hk#4�����g]ߞ�4�N��)sК���{�BǬ���ے2�d%�����C�d94�������a�#�E�ۈ�����)�P?LV��!�^vp	�W�����F]�2�ΝPH�{Ջ"������MM{��R����,��?:�t�����k�Y�lم�0��-���'�����>�Pq�Yi5x��4!+�#�S�~H�1���%@2�3�� ԡ%����9��$�� �d����L��8���M�v��s���5b��KՕH���{tӖgN���Ⱥ?��n�yG�&���l�D',-����sY�(溑K����?���48�L��7�\8:cE����5��$����H]XP�W�����_0�i��;(6�6�9�� �ԍ���L :��t^5*!��Ϝ�@&�\����v�B1����p�_�1�,����"���(D˝=8
��E����D�4<G%�\�¦���2�I\¹c{Y�{�n˶ ���ς��H�2���?�۩t�ɗ\�^|s>v�m����隁��%A%V�L.�%�q=�eOl��bz+$wk���/g�^�xBG��ĸ��!E�v����;�p=�cvʢ���>_�*�F��s�k9���ڎS�S_�6�gb�^�/��gב�1�!�[��-S�C廅��7d{]���2��t|��hR���K���A��)�k��q�P���J� H����d�fp�e7N�f��K�	5�8.+���KQ2g��_Uh��V�>$/���<�>�-k[�rWp���3W���r�Y��8j�#�yv\�H'��&8j��-�WjtāMf��a�*(��A�+!Y���.��aϢ��J *(�.D���A����D�w��`�zp�,w�,,wkR���ˢ�`Xg��_)W�
hp��ܳj��5+�T�[���lnLЛ��t�)5u�Nn�+샛H$�c���pis�j��<�뻋Z`#�(?c�G�UxL���
0|��EW�</��?S��a�_��֠�z��v0e/W �px�L��t8��2����`8����+�R��K���02�����~:�37�q/&!����2�Z��=}Z*��B@C��-����yu��B&C!�V%a�O�\�L�a/�"�%���S�Z@sd}4]ƾ$&5�8��7 y��0�2�]wY�<d']���J�ӊ!A�*�X��l^��oԪ��G<�F+�)��{}����]H>[ܫ�@�E��赨M��-��k��ɼZ&#�]e+OOQ��8���E�Pz;*W��mW��"Zҟ�5���!C��t#�q��p��cKtM\pqh�్J	� h�\�DY�Ca �~�U���L���O�žNJ��,�іC�71����̻���Sv�K�.H���6��0nv�j�:h�����g��)��ܖ�Y�ˬ��7�n�z����y��m���z��6e�S5��9��]���߶$ ��x�ǝ9�M�^fB.au��Q�V�ϩ8<2ja!ԵR��kP�{�7[�m�f
:�\T�@t�/��&���cn�e�����VoHT�=��l]&�.��^Ǖ+|��U�4��`�����
z�@gp8#v�W�<(������*����o�A�x�U U��:���Ǳ���@���Z��0��=Gg��Qv���f����H*\��U�@JG�:x�A/�%Jؘ,p�J����{$���G��	�&���~��a.�_[�o�uo�A���epW���N<~o)�H���.�`T���Xm��ߋ�k������{�/Գ.y�Z���S���
#��vZ��ky�"�bO�Q�ӖЍ�j�$"8a�X�KGh�A��hJ����p/��wI�!Zt'�-�9u���Ą��9䂤�ȁB��t0��Y:�{f� ���F|#��ew)q���\���|b�i�1����g�Ge{�����<	3��u�Ᵽ{������"b��N��9��7W���K5���8kQ�<_t2���'iAW��Ћ���,��o}䎏�Z��3b2�
���8L�
F|ص��u��_�.�EG�$]{�[�Y
j��Q����3zB��N��.b����my�z�r[c_v�堺8��c��"brea��kX'�E��ہ��l���*�X�$Kw�߁ '�j���==tCs
:��Z^4�*oĕN|A�?����q��!}Y*��}P�XNI����&n��4�D��E�L-�_���3��|ծ�z��y����H��R�L|�����af����N�� �1�G=����oʜ��N���tߕ��_��Qu��c��G7pL�AJ��kn�\��h*�`�(� ���Ư��mkUl�r�m�
�( �?���`m!Po˭M=�D�pStmTw	o�ǩv��w�B�����{k�,� �oW�`ΰ���`�k��AY����t���'�=�P�e/���	�+�6j�p�^��.�]L�v�����P��,S�M��5-
����]�MCf�����g��8���[�ӢUn'�$����'�������Q��(3m�b?��0��	�Q���η��X痆>fV�Գż��p�$2��훾�8�A!�-��Us�8E.7�]��6�,��P�<T�k*�=?�T|��T0K~I@������pX��N��H?�4��k�=��U(����Xt������_7�'vSs��$O�	����9�����P�G���2�c�E&}}�l�� �nH��sH��u�J�L|�l��-L�<KL���>u�x&���U����ͤ�UB�ˣk��u�׶�p 1{xߏ,��$Nu�9�\���Ŀ�R�����
`O)���wϘ$�I�]��a���n/9y\*��)Y|!���f:��8.�~J���x�ϲ@���p0��T���1@����Fu~��b��>�V�t��&�jS�WQ�b&]���F� L<��g�k�-�lQ�$O�	�(A��̓u�h�����
}qk���x�0����j�	{A<ͨ�|�=\2�ɐ��������;�\)��_�'9�Px���&��ѿ����Ex`��B��La�L�S�M�`���!'��a�����0���Пf��E��F��z�Qwv]�G�ecǻ��>gu������F�:Rf��5��f�L3MC�<Nt�C��!��t<�Y!��R;];�Y����^t[߭B^S�����i��]��H<ٞ�z����8��0~�!�%'��bpC7_a�Q�ٌ����i�^�ڡ'���^�dYQ{S"<q_]�+e-�%${����B��`G8
 ����6���%	�,Q�{22��jW����H�G�b^���s�HR��ȼG���x��2�q�Lft{5�>z݉�u��Ĵ�f���@&w�±V��L���ʂ�����&����zfo`�Z1���\�Y����V�Z���'}�|ţ���}k��Si�
�?s�,�ADN)����ʮ�������K4�0oa2��;sڥ3�.GWY��LF辋{҅�T1��5�.Y�gWRz8J'i_ק�3�w�
�X��e����a{��!k��Hz�q8.�m� Yﺡ�_�N:�֕е�'y |F~
2�0@��x�g5��[}�A^�B�������vj��5�|��v_:�3=D�q�������/��_꺜���3�Vۦ� �!��-�^�	�7p#�	��6#x�Jc�qQ���jf1�5S$r��!jPX��g\k��r�n`tNÏ8E�ŰV�QH�c�����` ����j�f��wqW��-ؘq�D��2��;Z��2dY;�&���H	i̻�8�wo��L��j<$yf�|2-�e;Ӏl��I`�i�1����y�q婩D,k:��Xw4�6'o��7:)�:�����!��wX꾘�%�ԔJ��$�˂q/n���1	�Mk�K������XV�Q��P���_	�M�)u*�#�#<�R���`�T�s�{�&�ŭvI�n��0������:{rr`�U��N���
!�������]+(ʙ��
?.R��$iY� j�3+��')	��A
U6�[�e�"�q��b�8��W�B�}隊�V�W*�x�����:�Ln7t�����zΖ�ǁѰIM��׷~@��B�|Pf5��ڏ۝'-�:\�����T�=-Y��l%c���i���Y��w%��3������v{cFoy�O����
+'n�P �Z�=ɂV1Ǎq��2N�v�I)c��t�!R��� �����YZ,�8&ΐ����HG���ٮL��7��l�^��L����8�غ�K��G����w;w�<	���ty�F�>L���6��i�����5Q/։�W�T2���Ü�AD�M�PhM�?xz��NB�`(Xm"�� Lg��|X���]Q��|�_b�s5�#�����X�w���S�Ax���l�T�sC"�j�g��̃U�A��N���ӬW��Y]�Rb<����Um�wJ�zoYY���$�ϒEXoa�����0��+p��bJ���o�*٭�_�_����beu#�=y�"u��WY}�@6�,�G�,?\�q#���C�~GuKG�[����wHQ<͜w�;���G�K(ޖ���5	�7��3�c�����p�.eR-2��d�`=�
^g�W�&�}Ώg��l�z]�V/���N���蕎!�ݦo�L�^"��B�����^��k=M�V9��R���ANrE|�'=f7����Bom�w�C�c�WI�h���,^X���l<F�.*N��e�������D��*�&��5][UE���W�u�E@f�˔8o�ȩ[��K��
F��QXJ�$)�5N���Y��N����O��8�r�#/��g��,F�T���/�R�>���֪����*�^��R_ w�Z���u�F��FI���-��odT�l�����Oښ�7��M���E��n�d�d@��A7&�C	�A큋6�ZM�Ō�`W�QC}��$�y(�xҶy��6�� �u��@�.��a�j+�7�\�:ַDg��_n��h�ų�8���	��i�wHh���^$%�8���s�W�S������M|��W�k��[Q�֨�W"�UAv��}�%$���:��茍+���i�6��nqo�_0b��V�$W� P��F���ͼ����A�Ў{�ژ�MQ���)�;M��F�������)
���R,� ������bJ\���.sd:�YP�0nA4*��ڝp0�����Q3R�H���f�/i���o��&nB*0��3+�i��-�'��/�>�/E�����{O�3����q�g��Ej�#�r�y����Fd��w�0�%}6�7r���)f���`��m+�1$�}��i�6��E6���o�T�Z�2�O$v�<a�#|�2��`OHN���푂���6��;t�ۧ�A������jh-/r�����l�6.�w~8"�/�&�g/�%�a�G�Tj�@�ƜdK]�n�O������k�{�]Y�Kы���:�R�����pD�v?{���_�qаOU���W ʵ�+ˊȹM�/:��H��}=R��� Ͻ�~6����MG��-��:�>p1J��?yq���p�9��ȼ�]�u�����W[.�Rb��@��Kw����E6�V-4��AcJ�f6X�������6��R�~<��(�+�2v�&+��(B�y��t�����W߷h`���I�4hߔB�i�HTx
|��ٓ��1uD<�fP�*I��w��L���;��PY)�f��%R��:�zK�L��h�������l��9e���u�e �S3I��-	�^)��Evn�9|z	<Ű�L�=Mp:�^�Z#g2�Yk�԰`��'��:��k7�v��C\O��Hn�U�89��QZIw4����<pc�¤����|��Z��S\J ���w����-`(�q`��C�L�c��q��L���=�ЃpvC�_�·X�5�.8�ѻ �����Ґ<��QⰼD��u�I��^�'M��}�z�_��f�J�������h��o�l��Q������I�3�9p
��?��sC<����/]Fl�}��B'�L�'��m������kk������d�^�
{6׉�+��4�+͊D	WhDf\>��/�͂,%��� �mD�Ǟ�x]m����yH�6��6�4�D��p�xl�2�ʴJ'��_�Z_%�"(�Uq��5�11�6�E *�Q,{3��'h�H���|��^%��X�󭧫�8�d[�e԰�Nx[��F"��s
��RI�"wM[�����lu�$�Ф��]K6jF��~$���u�
��{���n��U"K�)o��p�<�F�n��&og���z~YY������bk��䞡b�K��W�Q�g;�Y6���������倲$n����N1�:�u�	(�d���V��h�o%KAB�H���0R��`+�0��d4�u�z�3��=�U�˕�ྙ�M�ϊM��p��~ܣ�Ö�~��օ�͹Ʃ�{��-|�+��jט6��:Pl5��9��.�쵶ߠ�Y��$i#�O��)��\w�<�b"HX�~�Nκ����R�̍�6�jc�`"�9ވ���HVL�vyt�}1���CQL�V���z�q<��/*@��V�K��C������{�d�;����z���B��{��<��w��<u�2M�T�˓�pחq�@_���Y��t����{:��;#I?��P�r��z5#���p����/�MoC"u멞�0��.I����"��!JMv�@v=}��4�5�����y�|bjd�!O�Y�C(��%7�֧�P�.{���ݢ�d���rq�Hx�\����C�N_�S��K$0�zT�����~���J�6cL�%_��V�6{z-�2Y"jL!�0֟\?yt�Wn@�H��lK8�ݡ)��t�ɮ�^��7h������F2[�n��6Ă���ʉu' K�$���/�lM[�=��g��u=O�<䅁k.�1�d�h�Ct���1�9����n1�Qd��A�n��h�]��[I�ǂX
��޿�AFa;�����ع�72�Mkg������!^��[��r������1f���T Ik��\NF1��'�N���zKX5�h�, �p��VZNf�Q6���>}����t�Ba3x�B�M��T[�kL/�!�,~#H�X�E�]�Q�&� %M�`/(aա�(��쾌IǱ�5�Qn<c:��ra4�g4"<��(�6CiWJ���'�O�+�{��6 H�l1BV�y>��,�!� �v�5��l�9��@2�װ�#����N��5��e/�z�l�,]:)0��S�U�1�ש��dr<�^�K ��mןkpWq�O�������( ���amr'ۉx@Jl)x2g?)�J�ۏU����ێQuXQ�Q�����«f��S����Au�-p��+ږ?h����(���S�U�!�#̓#�q�#�tw����q�pN�tT1�p����E?ruL�h�*��
����Ŕt��>hV�>W����ͼ�����4��2�.��t{k����_wJw>F��������M���]��]�0��^{i�B��uUE%��%k�W*��K%!�x��
@��רGo*��1��逴Q^	�I
�#ӻ��@�k��#+�ʛ���$-G���d[dO�G;4�ۗ��� ���z �k��a���j(.@୤�D���c�A�kk��8��0]����fJ��]�6UWU7h�j�����xe�EWQ��m��p=\W4Q�@JW 6`|E��|�><�T��R��^Xv��|��aYy�{��7��y��J�y3�ur�"�r��ncqX���sV@5=�)i���^�Gͼ�,Ld����R��v��r�>�6�n�uL�4Ϲ����|,�*�b�mQ
c8�T/�[�V8v ��H~�u�ea�3|�9�@��}�M����7Eq?`�Ǆk�bl�}͙#�+zZ�wN�T�E)����n�=�?g?��g��I�%G����֍�!쌰���!#�,g�O�i���##�2����Ų�W����y:𷄦����*��M,hN�L���>`	�J�;b�G���@
����k��Ҋ^a5�4�H2��7���@k{Q�M�h���M��V��i��p�ز�w�e��
XS�˵��x���?U�f$�$s���^�C��S�^{�S�b�K1|0�\;��c�� �r3��s��
>8>�j0�Hk�>�#�+
�c� V�}�B�� K�O�o��u71AY>h�6R�d8'���GnS�c��q�V��3b��Mχ��,���iPʱX.����:I�4}a"��rB�j�P�=�h�Dז���f�Kq\5G�YVV-���L�ê{+t��i��U��M(���om%L֪\ �t�h�
7KR[�͎��p��p>B�	�8lͲ�'�ֻU��0V�K��yiӷl2���s���b���xt��Z�$��r�$П�Ĕ55�T�Y�&'�'�ANn��<d��4��Cچ`z<
�ؤy�p�]!i�K1&�>�,�8<��h��;κ��n�{����T/1�U�������_�5+����A�m(OS�=�d��%��A�� ��W6Zwt0]�����i�h�CG��Ǌ[����Q0���qx������5jS�a��Z��Z?�^X�ɱ�!�}��
�ח>=�V��v�]��&��L�w\���F_,��*U�C	�f��J�X�<n������zd֤����#��<�=7}��{1`�����Ď�ATr�&�aH�C5e� ƛ��8m'd��$�@��qɍ6it���7(���U4��N����{�s5����Qu�0 ����@��"��iTz}i�Dо�#�B})&l b�	�qn:u��P2Q��vR��儑����{�-k巰J*Y�t���d2A5}5������Kq�+�L����^9�3�P;���� I�ċ�W���N&�8��6>���D�A�%��I�B�?�Jz���h��,ӕc��QV|Ʊ	j��#,�����"�d�ʤ#�B���W�3U�[)�IF�B�0F=��>�}���/:js2�9��bV����<ƽ8	�`E�]  �a!�G'�~i���[�gPҒ����ִ*$���k�j]g$Iʍ��Vyx���� �/ǼK�ꨋ�ʣsӝY�Y~�i�T��&�ŏ�IN�fwf�Iqb�',"�{q(�Rl���h��5�G����{�8j��t��%9�J<~˙v���*�^ҽ�Q��geV� L)�䮼9��� �Uj�]�O6�nT9��AP�T�iI�3\�V�M���ބ�SsWCf�{�*��=3�bR�(z�������$O���>J��d�y(�<��4aM����c'z6>OS�BP��r�9�"�LG��'�g�Q��\�Q��Gl�|�����7��t��e�|Ť���5���4i5d.��"|R��ŉ�HA9˥��+	L�e�#��WEZV�t�l%�;���N�!lJIK�Pa����,'NKDJ�(��.7!T_�ҪK�%�V��ȹ͟b�{_�vƈU��c��PJ��"MI�,ܟ��qp0��4��|'R-���˛!���B���Ý�4�͔j�<ļV3�5�/�%��ɵ����'�M�J�!��(x	i��l?���A]��mK[K��T9&�1u�Ņ���>R��)£�+6(U����Γ����>��n}��e/��^��������')�,;�T��P�ǚ3��M���������\�u�C1�������Eݲ�k|KW��⣨�͚����)�-�_�]�v\����\:7����x�?)�[�"V.pV[nk�g�E�rq�6�koaj�t�D�D���<�@ 	N��Q���尣��LuV�G�U��������46�`Yy�H��gJ�>�c�'�؞�Y�Q5�TPI��n"{�"T�3V�r�5,M��Κ�5ґ{C�9W�$��ǃ���%X��ԓa��U�)�t�����a�\ρ�B��B���6��p�g?�]7$D�*Q�T��V1R����q�5�s^�)�_ټ(�H�e�}>���('W��%d������X�݊w���lES��_�	�x�*��jM�C20�ΎI����	?/�$9g�rS���ƭL�G� �s%g�r��W�	�z����#|<��γ� ����&S	̠��t+�.�;i��$MQ��&3��2���(ٔ5F5p*��*�7�/��_3o1J��rH����ɖn��+X���t�}<��~�dYs�̃`va	6�譵_Һ���aH�]��k��LT�$���E����.������}��[��_�m�v^���U�������T��9#�C�T�B9o^��|N-SC��VQ����߃�ꎽȅ4���H~!޺�2�����S�)��T���D9�eT��j�W2�;����Zh|���^Υ*��J��4�;D_�r���~6��6۔���pY��欪�,Qp��6����QN	��A�{�!:�����D��I��r'J�\�r�Qd/S'|T��"(�S�Ȧ&�q�}5�Vt���g!�t�'�c8'5�K�"pĳb)`ϊ%%H5����
;>'��2�Dŧ]��a�7:�.���O0Hl�5��&E�
p�I<�[�+���:���T�"kA]��43,M:뤤�K��f�Ui҇}�:�PrC���l̘���T�?�?���T,�i�4���`��L�����8Nd�\;W���|� �P��C������L݊��=��U2�{�Cw�<�g�1��N}����J�����`9�r��m8S�{R$>��8B��-�@�썞��3	 ���*�|ٸ�B���OEPP�M�x���Q(��_�D�2S��<���w�����U�e�B�i����-{���їF-�"iD��iQ��a}S�W_<Kf,O� �$��9Y|+R8"D�Ȑ=4
����
ȍPľ'�B��y��j�vI/����b�<;ÐːЄ�[ eQT��T`y���iL��{K�'z���Ƀ�=�Q�׾���w?��nŏ��;�㟃.t�XuB�T'�Jɏ� - H�u��_��6�IBP~�~|Sj]L,@�� �����qxႊz�Ge�+�1��+��8����>V��8��G�H�31	)����tv}mK�M��J�k�C��+�Lܩ:D9Ϲ���2�Jb�b����,WAע��r�j5����X �X��΅���܂���r���^K[4��ŗ_�����Fކ�~n+	�m3���%�	�®���V��ǹ���8����ٜ��r^q��6c��G��ۄ�%Q��hV�vLR��x`9���|��yt$,3pV�r&	�^*/��r>ٜ�?�3-��o2b���5�C/�|Uj�b5�κNy��{�u>��vo�	Yed7��j.�\�(d���2U|�������6ٮ�S/S$I���
!���:�o@��d������nL�pi�|^J�u
j�_W��݈*��,D��-_$#}o�X���kTy��iMύ���a&H)ͥ�D�A�2�F���#�wYb���$�)�7���� #B�<1��'�/�߂}=��3�N"U��1�LP�y��dIc�vao/)����ʂ�N�;��\�����)
� >o�}���������%R
$��Y�n���o�̛����	Z����h��8��QW�O0q��tG��@ap@�;R^b��T����'z��r`�#U=<���'��T�VU8�=��mhS"���/�v��v�U�������w1��4�}�
ւ�@��L3�6,�0�bZ�E��ѯLP����T���*b�\���!B-P��t�#��q�[��H}.���˔�bRB=�H��_���j��0��Xs��1�ђM-O��Sy�q;�[J�}��dj��F#������>����g`�p֭��-�z�_5���_�=���C�6X]��-a�W
� Dk�l�>���d�q �3R.�p	?ݻ"���)�"��b��SHt�� ��d{?��xV����� �w=]��Q/H]��"}�x��l�}'��b8� �� P�Ƒj&%4W��Xz�[k���UႷ�N���0ב�����2�O��̤!j��M�v"� ��!hHv�]��\�������REyyX��<n3j�6|i`o(D>!���p*���Nu��w�#i�gn�c΢!S����5��Irnf����5:Y�z��x؛�{W�x73v�ٛ0=�6u��@��Vl��B	[g�ϡY�E��	r?�X�q���ٖ����wx`��0�k�Vv���ؑ�rGF죿�f�}Y���!9��~=������
�+
��C]��@L�P�!P�B?Lz�9U��CR�r��]3M5?��z�Bf1Ob��"8�-S+۝���{I����Om�A^�{Ȼ�0iw!�=!�)�����ua7۱���t#c\\Q�GU8�\�m����2��<����.��G��P�lH	�`W����&�o�=�=��y���4�X�r�=����N��@��Z�;��U�ШH16�q��Ag>V{u;m ���e�B2��x��$�Y�� 3_7���C �J�Oy+�Z	��*S(uMxw
;AɃ}d9���Kꐧ��T5���������bs��_��w�F�.k�z�����jW��1d�"7ǌ�f�����_
�[�לR*����y`̖�i�1��������^2������K{�,@P��PUZuk�H���q�f|�f��.q���:0��@���X�Gm�����_���[��� ̎���q
c�����N�4.�*g�uW���v���e!	%�(P����h|��r��w�D�H:��c�yH��fG�rl$�U<H�?�6�V�M�����,��g�Bx����1[�(�Q����e�C��3a��Cm���JC���,�����՛20�!�E�������B7J�.��:§�o���Vo��0d������/Yn���T-e��
^�N���FB�2I) ���r.�X[4Qz������/{oA=�)u�F$�Ɓ��M@s���*��<-�J��G�k����%��yʉB���ëwbYe��8j� �	 ���_�� w �`�suN�� �`ȕ8iq@�D�9Q��F�;Tޗ��_V���g%-�CB@�nu�6�	f���h��a3 "�t���c՞%Zz�;��/��y�D]l����$YI���I��#�`v�����O�#��r6��Te��9y'��$����<�4z�/���w:��*��MXE�0����;�O��e���F],��x�o�r��k�BʙS�<e@�O�N`P����;7$���evpJe���r�{V7Q�9+�nY�t��I~���}����>��u�-\�):=����q��l<�F��|���GX��K,�c���A�=��N���@���ˮ�fF�[�M���`����������>��v�ʁ��%[�綊[Z�ugS"�����]��{�N¶�Ca��O�h�E���h`�u��7VToگm~L�a:�����ڀ��;��/�����vM6���(œ��lI/18�}D`�ľ��QS[�d��6$����� �
�M��f0�Ѵ>����w��["�TkF|��^����{P3��CR39�?U-����Y�iX? ���?vɗؙ����&3��'�LC7L!���ǟ�$P2��.��M�(� >��-�/3���A[���3�o�AI8�.�i�Ɂ1ث:
u��C-���\h��Ht����v�3���1B�o��ȶħ�W�>���ᓑ_Ӷ�b��V;�.�V��U�G���3�	'�g��f�:��ڢ��� 0lTۏ}�=�R[�%T����,�?�~���˛h�����xQv�N���qB�5$�m��;̳B0����}J�k_��l�=�*!:��q����χ�A�?�TЉK�<R���3�s��RKҍCms��2W��b�ą�˙��
szDs�43��m�W�7��]C@ s T��v�� {��Q�~�K�MPD^������t�}�°hE� �m�����E$[�F>�=�X�d���K��/I\��Yח��(֞�a��Y���}�2vZ��� �����u�k��ʞ��:���B x�'xCcJp��h|����n��}Z�����:h:�jB�1w����TB�7�h%�譥pXղ�7� �S*>8F�l;����(�Պ�����
/���Û՜�Y$Aeɠ\��+�������=�����O
�t�&�u4�͋[�G�A���3�X�BB-O�W�]�՜O�8�hb2r�e�YMOM�c���̲�V�˅�L��c�b�]N4e k�/�u-50�l�ji��ާ�ۥ�2j����p��3�Z�M{G�yfSy���#97m���`�UxJ�Y�T�����k*p���+�B��M�=�lb<�b/E\�<��uQ�ZFz��������'Tv��9�,f���&�2����������^K���H�Su�Q�N�(/������z9�Pl���g��D��j�P��\�|U;���wC���t�lCh��$�5�~�M_Cx������w˂�13v-��U3~e�xɞ^��,؝+J�sY�Bh ��]U�= �[bۈS�%X�i��~r� �9��G�
AyY>���W�ğ�J���}
DF��,K��#������Z�H�%��[�X?��˞ɷ��Y�ݢ'��`�0��ʘu1�����9���	�r,��r$b�y�`Y{�����u~?�զZ}���ǲ�t�Q.n<�v艠h�6<W-Tg��lp!��+��F�?:b��ts`�ݘ��U�l?��
����I���8ˀ�H���j7c\hS�� �R�m��@z�c�[�o	[������M0
�\�5�#��z�S�h���L��-�a,�����%��l��Y�fȤouq��E���r[x>� VU�\� ?Ä͋N֓6ng<�v�ۯ�, ���ra��e7֕�G��|���u�Y}
�M�v��x!����!,B��p[G���l�W(�����-da�%e�D=��6Ã�+��n�
�[f�)jy}ӓ6�x�\��:B'k0.�dJ��o$�<!?&PA��m�c�N����h EKǱ@���dr�z��ipB���b*��T�^:YlDNι��Z���^~��ꉼ���`&���e'	�K��V�s�3Ǩ5����+&Q:���]:�C�	/#.��{o�d�1�J�t��@(�k�=X���H�$���'�./����نj/)V�V�EU֎&=��B��NJΫ��J��N�G"	��c�5�����0w�~Ħ᱊C�B�o��%o�.��'���,Dy������I���+Xg�/��sqv,`/|��JfYf)���6�2P�����,��^d[�v����̙�?�*�qE�
����çU�W�s`�������#�y���eK<�t� T�66`T�e�r��$�C��-xV�=$����羯Y@��@�M���k¶�*.v(���X���B���k�E<~�	�h�������������V�ӿ
�δ3@���yr���6�k9Ȓx��M���_҃��#��~�9�t}����:�V7j��O��'H#@���Bݙ�2]� u� ����w��R��CھH������+#��P/�4!(ͩQ!y;�S3]�/r�[?~�=-��Α�.�{0⃋(�ɳT
���Ґ\�3�i���EGii%��{��{/����n��]V�v���+��U>,�:�q��W3i�Yl?0��JA�Htf�l���(�c>�mb<�!�2�(d�r�M�u�a��t���!ǋ��j j�/�@ܴ���6�^`9�+L���m/[�K�ڦ�f��ܧd�������N���O1�S�zE>�q���ή�Ű�D9D/�H�D�ǒ]���r���\���tp�v����I堝i#�LHg���y#��~rv��i��m���AA� ��ӚA9�و���JN�5��?�؎�_�ʅ,�ܗ�Ώ �0y���߅�T<�O% 6!w�h&�ӝ�+�s~ցͮ��ș������l3�%ؘVy����9�Ϗ���q;ʇ�擔P{��~;�M���5Z�X5��(�Z��{��.�HWw�����B;?�J�ή<)Fri�W݄S���+
�$n%��g����<�j�Ouj�}�'*��}j�~������p����峦3i�#�LOy��/�͑�9*O.|DCI�@�9Q�I��(`��<1��չ�qCW�������kl9{<���W���µ\�%G�{ٴ�@w�NYQҙm��T%��ϊ	��ܘ�M�������PC�.B?|r�/R��s�{�zen��� �򱮵/��fBFk���]�܆M�;��&33��o���j\O���8yŅ�.Ƞ8��|wX F���=�!NJ�%h���PP+�t�:g��IpM����LsK�o�#P��`���N���2(\���͠���N�z o,���X_';��ɸ4� ��Vm�@��&�I�dX&�â��A����ԧ僗����
4��52kF�>�>K�����W��4�ac3:�!��wp.>[N��^�h:_=C����ӞK�;��a�X����d�dx�1�$4B���c[�Q�_���(3Gn `V�8�X2!MK��S���Z5��`X�QLO*��]���
�q�nj�J.ɹ��p%!�H���JDm+��(ff��d���.ϐ,�V�'�)_����6�.��Dk$�?����ۅ�	��W��ޭ���;:̔$22[vjx�=f1Ƨ:�}3�m��]�,��ݣ�:�[�c�pO}a�l��_�~x�_dv�{Q�. ���c�Q$a��H`���|�_���R>f~rz���q99z,��S��	�p
��S��,�����i �;�4���Ce�FUy�Z�	�g����cdI�6��>Y�؆�_T�4VW@�3������ӗ`� ���z��4�[�����H:,��sY�����d?[�W}7�e�Fڷ,O���qB	b��R�÷�kJ�U��%�����y��M/��·�Z�yu6!1:��B��&Z�Bi��fƐ>�#d�M�GN��"k�y�C�:��v����P�.�c6\��J�rвp��/v�]�P\4.��ˀ�|-��)V�͹4�G�����~/�ކ'Ll;y��(�݅T�Sgl�I~|ݲ���w au�O�vezM��f��42c6��D�[��a�}�Q }RϠ��[,(�|�Z�끁SF ��T�V����X�T���7��W<����s8q�'�始,�<��}f(D涫t\��V��fI��^@o� ���.J�m�Y��<
����\����l@�V�+1����Ǭ�YQ<�2U@9i�սس�l�_�p p{L�2a�݂���05{��d~`�B�X�t �1�����i���f�]ȓS)	V��Yպ��@)�U^�W9�9��
3���y�ƩI����^��M���ʮ?�L������Z��$uP���K�24��P��y+��Ҿ$��f���).�R�&*���FP�P]�S��`�t��!7
�R���2$]�E�[�T���m��e/�U�H�g�;b��'xa;@�R֣�)o�0k��'n>�^�H��c���3c�4�m˿��_&x�6���\)y��t���R)߁�1�>"�B��y�j���d6 <�te�o��hJ��aWt��gwP���7G����:T{m���Kq�e1�b�<u�NQk��EB���̱�5���Lh
��R�*���Ǔ�p�7������+�{sK[y�N�O�R�5Rxd�oBE�(}�G	]ǋ�[���۱�R`e�g�{����75g{I��eㅅ��繾��%�xF�}��l��+Vȿ���o%���5��U���8��o�,��k!8;�S4� lIp�F摓�E"?��8�ђ*V�Pl4'ϋ���I=Az*�Xo�=5��""7�s�^��d�т$���b;H�j}�z�.�Ր;6��!
��T�9�g��t1�b�ucdBQ%v㇚��D�y7�%	"�@E$	^R�<�pY�F�!����=p�[� ��iRd���1�84{�gN�5�fSA=�~� �$�NRSj�O��5{5Z-�%|��8����(���&���I*�T	Tpӹb���V�L����d.�V��[�ՏYdOe�������0��UJٽX��=�Zrm�"%�����]��_�$���y��*�,%78�lSx�"�)pJ�>V�?��Ĩ�[2����߰��҆X��Ѹj`,5|���O���H3�Jpzh"I�L�� V��o�|J��(�ps�IFN&��u�B���7��{2'�7��u���^��'
�pXơY�C�`��[��{�%`y��̽|K��
��>��CI�m3��R�5َ<�R������Z��m\ox�ٽ��eI�ځ�5��D��c�d�S-e��u5P��(���kD�j���+�9��h�hv�����#����ѧ�I�
��O7�F����E�J�8�4h1#�xmG�����U|2D�](�op3�`��&��������l/�u�Kj,������Ǆ�h���(��6s mSfЫ�Y�a,��MIkI���=�?�����Q�w�����=ȩ��������s�^rܑ��s���n�
7:�ه�2AX�Sco��_�k[���C^���s�Vl�f���*����j����e�1~w���������/Q�5�74������<O���o�6�-�:��L		91e�E�q����>:R���}9����g"�f.�(�A߻���w2`	�˹��מbIK��k������������#R��u
<)Tz���KjާB��:���R�Q�i��oN�Ic!h}�XT?��,	k��,�Vԃ�i�$8��o�R����]
͈&p����,f�1��Y��	?�R�y��ƬG����hw�9_��M^ҝN���W:j�$�����΋����c.X�D��8�JW�nI-ХJ��>z�k@e�Ļ�����I�HcL��J��B��a� ��a?,G������_�ɛZ��P��?5}��hJ"d�g�:�|.��qs�����8�;�Z�j[Ӆ����g{���l�paq�X�:��F�����X��;C�^�o�G��F��4h�Bc�

� ���LL�.C����C�d�eFT�-uv�0�e�,���Ԍ02�j�BD'�?�����H�~%_D�.n����������[���<�U�F���2X�<
%D��l�	�h"�5��w�Ѹ�uN2lu�*ux����D�R�ƛ�J4 �U�"�I�ͯK�c��zW���1;tl�4�J*�;�&�#a���tf�0-�@��KY�@N?^ڳ���e$�J�^�|��۴���ht��^57=����%|�2X�ޙNF{���#I������J�Le�A>��$�ޚD�s�j��=�L�z~�>��wK=~DK�,�9;P;|�e���|�T���լ���N����Z�PҮ��qHw��N�w�ŧ���GkeS��L���*Pl��l�c���N����N���.�{P
w��̭��
`EZMŰ�/{�+��3d�^�i��?%+�a�نZd����@J�%���GCB�dx/��˾�c�T�l��LHB��֧47�~}_�y#0+�TR��e2���Vmi���~w����M�c������/0��X_ʼ�A�M7�m�PP�2�����TEz�X�+;*���� ���>�7�	�PJ˓ojl��WRÙ5M�@P��iǞ%���)��	�;��v���O���Ǚ�"�S�G����w�����x������]�Sb#N�9cy����6b[K%O5�e��}�(��yV'g�>H��4��.z���0t,�Rv�\>XE�P�̪�E�1�s"b�CS�8�`�af�Y���cVJ�W�{�|}���wOzQHc���=ߒV���4�A�=�Gn)쒰.�R�E����:=�G���%��D#��ɀaD��[B���ؚ$ƚ]I/�6AlR0��:Y-U?��ġeT�R���8�����m$=�@�>`�e�B������ʩ�ү�#�FF��xJ�������iDJ�޵���z˪I����]-O�o{������​,�	.}�8�.�J ֳ��a�U�(2zF$��ū�}_-7����{V��~B���e��z4)�����1��{:Wr�_�(x���&�hM�X�&�M��:�CK#2Fz��r���7\zHP��-���|aw-��(���â]�R�Ӕ�a&�go�&�E`�-���9Xv�t
�*�i�X�8NTP�H�VͶ��-m�	<{&v��$�Sg�.���S�A��i�V�2�~����z�7�1�;��D��l��z9��!����h�!0�V�O���(3��8�-xm#&K�?�v��L��A�(���u�l��+�i�昆9�WQ�6��*��2%�u�qN<�;���8�W!K�-bF%�Pl	�4�y��8�Q�s�����O%�Q�p+�3���|ݪ�(�A�AH��fj�P���H��"�{b�,��&k{�\��E��^�7�U��,�U��%lN@�u��i(pA�f�����ljE;�
�NQ��?'����;=K/��Y
�����r���ɦ�jO�>��(���O���^*��� I���7�	|���,L
HO�اVʇ����8T�П��1{V�S��m5�,��@�?'T�J������na}����-e*��ǎ����C9������Sҹ4�}И^8�Ш�st^@�H�R@#�b��:��y�����N}6A������C'�=���/�-�+�����u�V�d@�*�U�~_^2QYR��Q��h�����s\��v`�Y�/��]���̀tJ�r� -p�4�F�@>�vY'5�y]����!�G�nJӃ 
Nu�t�61��i��D8t����4��F�Q��#�<*�i��X�i�]������F@�� ZB���Q|�U}���1���UZB|�P���w�{y�r9e��%�����^$�+���,�?�)_�m��7yF��ᤤ�2��nGA����p`u7"|w!���fIg����=����1A�5��n~�_f�C���x�x���t����Gv`mY�����=o�7��&R�e I��Fl�I*���y[��+�r������x/�3)/2�u��>�O�M���%��!Z���mp_�s8M��(06B1�L�EliA[�#ާ�ﬧ5gBG�����y���0Z<l���A^X�+�,�Jb����f+��B��3d��XԶl��$�K�Y��F�����k��QW�<�I�����7�gDs�#���za}��	>�ϫ<���h!g`��֖�%�&�-��=��E�D���S��o����N�'��N~��<�@��G{0�q׷�sQ�ŋ��t�2@ >#������$r������<5GJ��qza��s�� �¸L�J�M��5�eGK�E}l��\���޳�ZrB;	ȩ[���5�c�b_t�T�n� ��,��PL�[)�^�
nNԮ8�<;>�߯����f��/7�J$�w��+d�o�2:��'�F�k�&�p�!��	�/c7ivESS6����A�-�#�����<��@�v��6}�O�a�X���	I��yK6~�}���߾<�z���)��,g���Ko�g�I	��aЁ��k��ـp���ĖB����(�����ޛ�f��W�Ú+����=K�1��1E�g�]���_�Em.M;ʔ��8"⦟P�OW���̵���*Z��M�*M4����މKQ!Lȋ�%�+g$>�� !C&��p��Z�_@ig�uf��wk����H&η�=�=��՜@�x��g����~U�lۦlW�/1V��P����G�44���1St���俬e�
��q��}����Ր�|׭��q :qǝ�v��-�ZoH&]n/�K�&���;�����D�2���-�w�u��C�칬x���Z�` R��*�W���䤋�P=�Ȼ8�����}�a�9� �i>�);�jz����8I�#U�_8�W��7U/�͝z卐���(s�e���0�m���r�OJ��/o��ݥp+*���y_*��)���0o25C&����Dy�
�&(�A$�JTiy�ꡪ*&*����`c�/)%�OF�����J��7;1ǵ��� b�}>^0��1LA�ͼ���}����;ίkv���q��Vi�ؗ/�zW��a\��zT֏�	� џ]����I�HD�Z���{X�w��,��ёCٵ��8�3	4��o���<l��|}��oD@
�mZ��+���h�YX�4G�Ė@IT�������s-uZLc�Fr���|K���4�-R�1�Jgi�V�42H[e	�h廋�n%�!���Й%�z�}x�~ ]��J��ߞ ��	��[*�=�
�G��'V�w�lV(�l�<"�b���~���,�E��A� ���b;��Ǭ��Vh�g�&����ݱ��c0=q�F~� g7�'䢓{u���J���r�r�Uf�bM�M��x�+�3b�j�ʭ���}^��&�փ�C?XXn�ե���8lY~��,	�q��v�4�"p���DD~��Y��k� Y�Q�&4>}N�1[o,�u�z��\���P�����hB��l��#$�p}1�Hm䉼6M_L|�s�B���a
"���@�b�'��b1�Hc>���
ۅ�XzPRߩȔ�H�6+�Y��n���K� ����;nJ�ћQ*�U;h�i_V�V��@�����$����ܥ38�B����ܡ���o��Q� $LY�+�Ҟ���		�Ve����h��!s9�Mav��]gd��B5<U\�j�N���@-BQ�-�m{'���3������D�+�u�����8>+ ���&z�m��e,��_�ӶYN��L��g'�4�oҏ
��U@��\HԜ8��E%SC������F�'�����&"^Y>AІ�M��M��ĵ�?[ջ�x[�G
C���<��P�W���������H-�������!}A�Bv�K�:݁���MG._�wL�-��c,{ght��c-a�\�`�����@��K�����  �O�4N����}��Lgӈj�0�UG��\M��CD?�SH+}��`픃<�4��ꆉ }���܁��l�Ԁ��#�cW^�'���ǐ�x��>Xҿ\��˭�, {r�3=�y��PK}��	o#�{)�Ez����uR�,��Mu���C�ڳ��"Zt�:��t9M"6���Lsg\�uN~	��n�F�ʎ!:Rދ�h�N�������?�I������RJt���m�va��č�hbg�,�˚^�0�p�J��^��SF��tH��F���)�(�d���������.,	�b�2����vd�1�( ���ӂ� �Dw��8��!�E����S�52ڨ^�1�$�>�{W6{�&x&nDbz�VС�+D0��,�KԱ��U�cF����A�V�;ٔ�,5�\��n����@'�G��	٫�G�s�E����D�(&;23�����ӗ�a:uK�үd4�n<l��*��ɉ��yh, ,�P���H`_�ԓ5���y�F/��ff�| �%ș���\?&(�k�2h���F|�ק$��~^�z�I����ܚ"���0���߂��*��TD�NahZ9A�$�w ��#�:`U���vy�BNR� �c����Ӛ_�uB[I�)�J��T�jdI�O>��R�Ŋ{�K�?W�\u��.�樁������?�����sĽ'�5��T�I�(��:�6���#¿tR�d�N����Hq�����m���,FO��Thc+�	��C��q�$(��"s��Y|l����̼�{X��f���h䟀Ws�jN�&�DF��Yj����"�5 �b�Pi��HO��Fv�7UR�g�T)�iN^�H���i��z��=9V��t��z�U��C�8��X*
c�!�8,�������m@l�=�/Ѽ�F7��������ϝM�b�ܨ����S޼-|-zN霢�	x�c$�����ZP �������;���
a).Q�*�d�:������;��+zN]R��(g�5�����r�%�d��V�c�~�T�J\K��f�g��?;ڳk�̭��T�?lh�jЃ�4���0���#�0�ǾT|��O]� & _g����������[��2�6�dl0p��M7gց�찆��H�i��_.�SXa$�[�C0��IֈG��Ga[��%/�U�r@�y���jӂl�Y�!�͂^BŮ��e�2��JP]����@�H���e1��\(�j��^U�ڞO_� �Þ���6'c~�i���Uȅ�y�?� /Wx/���tMl��	��e������]��qd$^���3Յ�����'l��;ីk��L�:��� p<aqwFa<U}�l���s�Wm �r�oứ	�����9���_�5�QX�ņN�x�sMj�Cs�ٛ� �}��/Ƞ� a��6ƴm����V"����C'��i*���)L[%��')�qgõMgYp|�D���K��%��92����|I�8t�4~�}w s�T���B�=RZ��b��Ok����h����B���M���a.4K�5N���wKB��<��R'����C����*����|�_�"����=�ݠr�����{�ue�����Y[��౤�)��<���sZD�/��̏!4A� �&o��e%3#�@iTtv"�{P�&��kəSZ��/��a/��%y�'b���U�mikP<0xFe�"aj�ƾ6����-V5;��N9��8��n���"����SȰ9�?g�{��c��@!��ǭ���y������G����K�g#��ouD(Q�~���Z�����@��-�i�����"��G�H7�<2�an��3���(�)�R�Ǚp�����R�jd[ -GÎ{�\T�Q��������8ˎ)����_�����n�ic�������I-�\H`#}�p�8Q>!����_��)Ó}9K>�]�.>��[��R.��F�hD*�)�.c�\� ��P�����o%+x5�6�3�oL���� �4Mx4Y��C��Yɝ��wA����s��ٽ���!�a\��W#�����8I��Ld拥"b_�P�gm~����zV=�J�����o�$�w�Sy����r�7��i�B7�-�`^F�Uݏ��pk��Vq�svV��Qe~�q��4���ؒ�#�c��L F�yYD��]���ι�7���d���Y�V�Ù�˅s��C =Ϣn]�J:���'z��{<��ĺE*�ƹ�����T�IQ�Y�#"~0�V_��{g,���/e1�]_ٖ9���
�j��_
v����,~�ڊC/1h	�f0*��%ɱj�����Nx�G�]��J��G��l8h7�m�mn�N5������cwg���7��&B%�Th��cN�� ���g-H�W9�񿼔LP�U!Si��O�[J�4E�h劘��n�
����^�
"���Tt�������7w���W4�ѫ���8�/3ر�?z���Z��1(�}�䈜�e�ֳ�T��Q]��>B<dh|�=y���Jhܣ{Wx�'���� �&s��#z:"S��Z��!�>�$W���AOz���m9��������˾��;bJ_��0:���Q`����'���M��I�/js�
W?�y�%�����TkB"��F6�R�S$� e6х�8���4��"��j���8�o����9mT��b���J4-�t��>��Y��n ��%�:g!~�"���X%�/>C:�bo%��?5
�Ϊ�)8�����oH�k�V�������5��TH�紦Ę�������|wi�%X8�S��E񃟵/�HK���֜`�r=$]$Z����AE��m��#���'�z��*�;A��YiUv�vE��o팷f�N�Bk��l�r[�^����YQ���)�'��4��n�չ��<+qphY|f�&M����5m A<���:�cȼ��������
}Y�"7���m��h�\��f`��!�<�+ ��!,���}��3�H�k��!+����A̫|�2�E)�N�kRj/o�!�U��񻷾ȥ���_�?�b��KP�M�.
�J�$��ln�-7�	fO0i��������u�@��tgP���s*.�(Y�U����&$��o5U�8����t�Wf�*L�y���O��X��ZRֶ�|;-3�"���#�]��g@��VCjkݩ���P,�m�<�Ai8�b�bT�TL��z5���+a�0�8Z�y_;���lSb~�Q1�� �����l=J2/����٭�-fM6�%9�	��@Ic�b�zL�����V�����Hq��.�3-�*m�y��"
kh1���/�\p�'���͟�a�D%
{���̬��aD��ԨF���j���K�l]:i���oT�tٮ=��fw]	����<m�w�&W����{����DI�����*�s�:fQ���nX1]Vfք�����V���T���i�Ϛ P��ߪ�,�q���=��R`�2��KQ�i���vNւ:#&&�߼�KЀ�Ʃ V��Bj"� �~UNU[C��Y�T�gT0���i����K��ا)��pN� 9�#^k���"8�����H;�b��?��c�rQ�xc�;9�*�r����Y������&�]qu*��?��"8���]�R�l,h�W��	�rJB}�0��pg�����:|G%��1�h[Ϳa�z(���?Fn�C��n���E��4�=>��DN�%���,ͱ�c��B�w���>�"����N-*��mx��q�.��+}����r����A�"U�Q�ԩOeE�_�]�W����ퟔ��E�)�O��ldE�~�	~��m )�[?2w�pt�j�L�[�R΃	��%���y�+pD7��@	&�`=�Vx�zs�s�m=8u}`8�z|t��=����M'7C]��
Ʀ���IJL2]�ŃW���궣�M�k�Vh��Dm��`��V R�`д�'^hD�8���]9�g�g��bm��^��`�i��ޘ��a/K�G5ԛ&�tn㙨7)9?���3 ���o�������3l��֓v��w�(c�Xd��	ڑ�sP�b�MQ��P
m �R5*��tH�o�G�Xaen�L�+ծC3GY��[hկ(t��ԙ]�R�?����ڔ�[ջW��ew¦Y�j�7r�4���B*4��t�������O�|{u�@��+�+�r�*i�zb�	2ES*�]��Q.�Y���C�T�T�AD�K�Oʍ6�o�L�85���]N���@dO#�L��5:���Pژ6�"���$��ic!;%�W
ÐF�@�� ���6p���ĸ��G��gy'5��9�1��t�s/i��|��$����Zn�2�x�����ly#�+ɶ7��=���qlyp��`5�M�����ex�^t6?cV��Z������<��J�e�\�4}[?�2	��N��|���H�{�w����ˢU��*6q��� �-��a���	��`ؿ�p��E:����ǹ�,�*�'�I�^U�]Sx� �^Ai	bj��d�������5=td+畊�sp-8���$�>��$b�Ya�C�[��]�����igX8�l�#��5���YoqPf���;�͢,7#��~�a�6�?�#����a_���i������ZHb0�a���s�;MR�������(Y�02�鱹%X�_A��&�A�3M��C�͈�˛��������wꉂSeN�GĦ�pD ��B���b�~lyi�����;� 5�B�jX�cy�5S4>4�9��Q��z��$�����Z&)4��m�@�&�Jm�Bq2R�^���������o�i�Nހ]�7,���<�n*�]- )��(GvU����9A2�̑J��CZ�aޟ2� )�	���9+Q�f�37-`���NvP�o�[���ud�-�'��o�U�V'��5�#�>��ӽ�?�-`�j���	���}���$��̳m�7#��\��bZ�C�c��pzY-#i�%�0���C�����gs.�-Cy����C��wC�:��fa(���jg�8�݂;a���� 3*~��P���3�*q�${iD�b��@�Jf�����7���5j��3f�}����Z��4Ky���d�t��7�i��9�	�n*p3I������z��%a��IT��/BՖA��3��0���, ���dyPMtA7~"����a�%��I&S�;o���x�P�B�����i:0.-](ꊐM�/���SMFZR[�@��^����1ѿ���q���%�`���"L^J]� ��L�CEn�o�[-�л�=��6����&�˴v7g�XEmZ��$sZ0<F��r6��kg쳪�R�m�d��Co7^��� �e,M��ƀ��]FT��Âr�7[GѺ�ͩ���F��?��*���%}�����+�D�I�Y�l\Ӆ��B�w���@�!X�|4=3*�Q54�{hgƝ�-��f�z�� �2�rYf��f�sM?�w$u�g ��^E�
U?���Ȥ�S��V�+/Nؑ2�N'7tȊ^�ƉDeW�VW��M�������o��e��"��J����zt��K{N	���gOM7iKP�c�y��������kԒ�ԡbj���x�:ݮ������Yk�߹����H0Q\-�����>r@�8��(��va�ԥ�zz6�ZQ({^���[Vb%��sPO�fdGӚ�i|�V�� ����_��`�՞���
�Z�GМ�g���rׁ�x��E۾���`r��9�M $[�0j!�C�p����q��nF����{o�Č�Nh6�$�
1j�%���Dl�״U��(�?�D����n�r�,G���vb��	�T�q#Ce��m�2�Ĕ�����;��2�΢yQ��8��O�[_A���yY�[~T	S�(u:�CV3/�OT��7���׶*vŢҟ�K����k�Z�u.=��@�������^a�É�Z5�K�ִ���6�Y2���{M����I��&��J�*:��1	��s���T�����R��c|]��d��tf����B�?�Zkd�<R�tp�z2��<�@1���Xe��?F�L濳�F���?�0e���8-޿u�m�;���@�6(A�W^���f
^nG�a�3��AГ�q���Hr��M�y-w���-��	�r'tZbPK�?��* ��o���@/�@��<�rHr�yD>b�f	-`�!�1�H�&ʌ߆k@�@�v���!;oG�
�m��04�n ���aou�w��8mҌ��p���T8_A�utG6}!-��Ce�3d��I��;�f~��Uy� ��	%x��{bz�f>�R���N�W����7��}݊K��!ö8�����rl��j���x�:ѿ�E�J	@\�Z	� ��)��=7>�Q���zk3���]=�72�tK�/�\X�ٙ�Ft�<c�ly+-|h�!Wf6� ε���u��a@�#S
�`=������JW�&'�V	��]XXRz���/����ӈ��>�$���
j�"J�U�f%��a�)�����	H��J��U���
��SX+�_Qz&�X�Q�s�����%�ALj+��у�9�a.��3#wI�s��մf�-�Pg�5	Dӎ'	#ɍ��� �?����6��=<�|`}�y�S����ԗ�ݥ���A��J=E@���Yj���8q�$m{��	�I����%SݴqU<v}�#.�<������cQ~��qZ��m+�w�!/��u�t�F������Y������\(�qW?%�����埆ƺ3L��P���"!Җ(���{�)��\q
	���2a_8���Y*`��4�8!0�Կҝ�����w���5/�Vs���q�y����m����2�E��gc����8�����@�"J���	���wYKg�&�(��?k����_��b ���Dx.[d;z���(kq��7ۃ����򠤜i���9���|Z&*����E�������J�|z2Yi-r�)���UVX�խ�;�q�f���ܟ诱����Cq��Vy����U���Z����0dp6�B�Y+Q7¥�:��{��p��v��nխ�"����]@;����N�F�K.�w
 ���P*�-����g�r��9nf
q`�q�|F�C)Q'�+��g>��ܖ[�v5��o��G�67�[�)��φ�V�a�
A�Hʟ��Ώ��l�[:jx��W[e/��V��v�6!긫YM(lJ|̆�7I p�PY���t���o�T�/�b�d���K<�v�gV�G��=���oP��[�Zw
�@4���g�	��A"��l"
)��W��yg�o��ה=D�h�p4��}�]�p���Q�}�:)��]V;�m�OV�s�	�Ƌ3n 04?��Wu-������$/��漏����P�{�x\4��0ږ�Mu���^A��P�����f�4݊�p�Y�M�SE�
>�k������Υq��U H���}���qW��T��[��K����5�i"vH���ll�F��!\�'�P�c��:���.6���|~���r�yG���1����+��E�lN�I���BUI"����h�)x���598��!�63��&��	ӡ���H}A-��4L�
�D��oD昩����`?=�BI��!��-���΁�W�y�ml1������Ѳ�� ދbe*��=���[Q~�k�����A�M�8���-��p��d���8���} ����u\���)I%�!u����ʹ��9b<<ܫp��.�PJSJ�t��
�E��:F�Ǹ�\��j�}��L)�e�ߒCd��m�+�O��k��Isi9��A
���Uor�y�O�3�G���4؇xo3�˴�4��Dw��X���r~���x�e� `̬֢�?H�vKU/���#9�������3Jn�s^֎wK�˭GK�ߊ�҃,���^��#CaU�J�[���i�Uw��[��ka�1�;Ai���E5�_a�uƳ��TuБ�BW�?痫~m1�d�qg���Q
QH�������ǽ��J�C@A�b��6{�#fY�=����������ԵC7�VN���1|�������l@D
m��-/��͠bH�#�v��S�ߘ���y^��%2�mD�مL��Y#��]jܕ��f�g��]�FE�ز�`ɟ)U\�!�,�o��c�W91j��1�^������ޔ�|}���'���?r."���ᆪ?�[�<u��ji�<�l�Y���P�^(���SE�3Hݿ��ҡ|o��UhN6�����>�qEN���҉>]���=2�s��9�;R~�"��'yB���ƒ��
�0j��n	�wg�6��A(�｣l?��ye/������6b��mfL����8l����a^�I+��#�l1G<iȂ�D]:�9�SF��	a��Qi�=�	>Z�;�}4�g�$BY���Ha1�/7
� �Q��$�'�E PU��	�bt�K��rp�ca�񫆶�O�����|kzhv���j��������R(����}�~JI�I�F�ۦ�G��H��X��6���p��_�U�a>�O �������[���a�F����%�\$�ڢ��j��R/�^I�{��>�~�s��s@h����&�6N�����z�3
��JP�%_��Z����if��r&��A%��.��8�WtN)͝�ݡ�"�ίRQ>��7~��n���#�O����7B��c�+;A+}S�$�Wx2�ٕ������Y�K��
��l��$m6��*s��x
��N��ӮTc���ͦ�����T��4z���w�.vћ z�/M��IH�L�];
N'xЂ9��Z'��C ���(�d�jKS~!�q�pɹ��#� /Zr5K<z�s���������(����hN���/֭���~�sq��;���Q�6Eu:�V��.lC��/:�j�����#->H��&�\zӼ�M� X(���\N�/4N��c�5�T����B�)�W�;�/ć�tL憁a[��P3�R��ځp�6����ba1+����'n�ȑ�Kx���G�P��J���t� �A�eÙ�ָ|�dM�����}s�R�:�R$e)�E��4[�Ƭ� ��_�@�������y���D��͹�䖶��l�
�A�ݠ��}ȽP��P�e��_{ �o��52����
5�ЪӍ'�"�"��ϸ��e�ʊ��^��8�3l)�e�|�.��\yWe��&�/qv?�5�,��5�E�C =��3J��D�|��ݱ�#"C�������bj��ա���r���g��y��-�l�����ō�6Y�7�������~S󥁂/=�Ö#��a�NH�W��V��C�(�-����%�o�hn���}�do`+���}�c���q��#h��f��Z���x[O���3}�V����H��;��7ʥDq2��t���R�
�h4²,��+#�r�`sӝ�7V��Y{���*���[}:5g�<=�M��Ȏ�y�`\��a�р��8��B_����[��f0돻��^�̼�no	�C��x���0`| Á��f�\Ka�dF]��G��+����e��}pl��Q���UV_��K� %��r)޵������않�@���K��ktԠ�غ���3�qG �aaEO�p'FL��H�"V�
�m���2p��71�n��Ʀ��� U5� ����uT�ٔt�hR�)�ķs���7��:<ej�)�������^#�rM����ì��ލЮ~M�_��"ˢ%<��+�Pu<�eJutYi*�+����G�Ϗ�O\��9�1��^���Y��/y����٣1`2ZԿ����4NGz��a5�̓�Y��f�)��T�z9w �Dm\N�q3���a^����`��D[ȁ\a��5�Jj�B_��U��Գ!��GK�h����j\\H���͵n�Ė@���f�D�4�^Si8
 �Bd��Ī/����X-\��AGj"A��GCKz���:Q�';�
M�D
���9wH�_�MSY�Rb-�i�_࿈ǒ�z�e�
��r��0[~ʴ��\��_�H*���e�LHn8�vz�v�"_����n�4��YME�ţ�]�GmO~'�w�2v�*���*yNt�|�D21y��&7��L�i���R���!���v�}G�H��e���@�M�m�?n�^�M~J�\����JQl����Y���.�f���K�u�L=�󵺈���~/,��n8������� #E���+T���6��d�l;YJ�吒_�Dqp��sT��r�u� ��k�����#`�Opܶ�N�3RPͥ&Y�qj��{���<n*5ج.��������.9]�?6EH���Z�ڡl�w"?
>J��e�V�eE��)	X������|�Ku��h�Z_UZ|��U��웻�}�uN�H�F���H"da��MN���h�L\PQ�0&�áAe
����p�Z�9
��]�I=/k|ib-7H�<զ� xy����
Ǻ�jJ T��-�j �%����Q���cCq��|��zf�X�BZ;e{J�(��3�{$���\L�Y<d>n��vZЕ~��F���?kU��2`5O3K�_����\��rT�� 31�
W�[r��-�3=8dH�,Ul4jȉ�Ez|e��������Ɗo�Zp~���95x$G�s XZfڿR�V�b+��Ƿ�\zu���˜��@ܷ��_#��C��ri%5�r�������<[9b�7�!�tb;0�In�%+l7X�����~�&���� �/�%l���j� $\�"�2�j��+�M�����	�]\�}���R�G �5�E���}��=�����PV0�� ��cX����}0�˗�+���f�J�H@�4<>8����E�C�Ӻ���Ė�Ð�_�G=p~�C#���G�>�8>Ǿc����o�b���?�\�j�pd����'VnZ�p�H�נ��������X�s4Du�j�GS[g'�br��mU���Cg��o\CƊ��>�G׹��ttc�Lc����F��,�N@��G�����o��Q"Zd�$��ob���v����C��Nu�kyP�����X�Cep!X��c�~��?e��T�,��w�=|��.@�;*�3%z�^艫I�	O�:�o�P��.��e�r��w�u���ɻ~�B0	X@��������Z4���e���3P+�M��$��l1�^��!"1c����KAŐX�dq����Bq]����v�uCtLq�m���T����P�إ�7C���Z�Y���.{YA�G�Vӛ�S�do7�S�>�B�)א�K���!F�	+��c�."y�F��Z#bh�D$�
I0�b�Sx�8:9�����#��Q�5%����^��K��y&�%u6T���'�� ��	'��m �p������ |��J�Խ�N
3p ���+�U�H�@��E�5�xÕb�j�i���L8vK�͘l�F���Z�32d�\8�z�L%;��흕�ka�U*�-0�"����9"�˖�n_]d]J���M��C�H!lc:�Z�<U1�)Z
���K��tF�G�����%=�����;2
%Y�.9��qө͝�[&�|��-��ˤ?'ef7|�����]`~"�Ö�<;д�@6�A)Q��®�C��)h��I/�,~GsMɑ��̓�U����ӕy� ,/Y���R��|��0�W�3�����|]kV�f���������H�vț�Z�䒴���~�aC�����1�<T;|���8��pa�)bo��Z��-�(�CZ�uF_j�3�̣����+%+�POVU\��< UMf���������, ]{g��?~��o�H�k�Wsr�j�k�P��I�è�z
�R��ך�<u�Ǟ�z�R����S8fn�O���)��ϴD�����%�����"�/��L�#�����{bv��|�WB�)��;�i9d�?���1�?x.��!�S|.�$��/���Y&�'���\䪂�������]K���E���/�H.;$�x(���+��=|��*�������8Ph�ۻ�~���:�DET*^�v�ҁ������������l"����/S��	�w�CH��cXMk6��7��%/D��0����9��~��FpXxEG �|��U���i�e ����I@ׄ�Ɠ�P[�<�r��|�����Y���o�2��:)�l/�\Ӆc����*�`'S��k�A ��Ԛm�>��$��H�5u�������!J��<��(�9�>n���f��Dۃ/=7$�vo#�\�/_!����;�Fx
#�E�'�Ė=��dy��bg�h:9S�?�:�W��ti�CĠ\�wj�>�����1͸u�d��
@�I=���������{+.#�����`�`��iF�B�\ʌ{�(i}E��VCJ��j�q ��Z�S=D��)%{4����pr��f��������E*�����	� �HP�d��J���ˡ;b�o[����E��X?��l����t��U�|W���[��r��4������]������M�yt2K�_iH\҅���6{�~ƿɺ�5H*���� �B���x���/%����d|��������r���d��ۥZ�s�z��,]E���w��i�Q�k���s�m
;7����ݵY�p�{�v��R�X����$�˦=|��l8.X
M�F��N��jU�w�p��RA��|��k���v��(��;>�n��3+��ń�1R�~�T����'s|����[_�Ț[]r�S���^��������w��+��4!�I�n�t��/�i~pڕ���C�.�W��p�.ʓ�������&��7}-�;�����R�'�{-|l����]wm���_/O])��m�3�����q���7����VG��l�v���,���b���5>am"��5�`���B�&��}^�/RE[�z+(@�n� �U`M���b3&g�0�-���j���F�����P�|=}��=�;Y�*v�rU�A�r��2I�)^Zۦ�	��aXd�>Y��@c�j�I���dp��ӴU
�#�o�f��\�.z�"�w��Ì����쇴%��ҝ��v+��fP+��ᬍJ�[\� �����f��RZ���|:��}Y��)A���U&k��;6�h�����ƺ~J��#����&��Xb)�T��vM8�]�H��8\�, �J)�2w7��L��'<ND�=�;m=+����2*�nھp0`F��U�neV�䩡���!P��lx\۪kA�-N��f�h:��&H`z�����_4���n*�ɩ���^߫�EJܝ��!�����[��ɖI'�մu�3��-��&d��yz�;��a[&����E6uX� I�'�:䗀z�ԧj#��L�#@�$��.�����H���'���O�6�(���B�wo���l	c}�������86�E��&��O�f�lfͭ�������x`�W�,]+2E�]f�%`6��W%YG �h.`sC�/l�yf�7��W�_���<E���/���4��óc&ƛt���:�9��3:�d�x�����3����rv~�ȝ�U:�}�g��C8��Q�!vYi�5�"uD��*�?ڦ�IdS/,���q2�m�B�B{��m�����������|ݽ�����?"�}����@����#�mõ��FMF��~̵Q���"N[#���T�������(��=�r��n�<��Pg�-Z�ư�1͊�妰�-��ɍ�?�Xr
�G�XO���s{���T��MZ����v��Ä�mvy��Ȓ?�(�t
��/�J���kE��K������Ɏ� �M\ݨ��L���f1&U���X�󵃯<yղ[7W��kj�W��J��&��V{$Q�o`��?ʇ[K�iDl�+��s���N�~�e�k�Ay��4i�^���u��!&4����ʐ3�Q�^�����W�}�0�2if���lC���;R_Kם�CE&�>Ƒk�3YSj(����s;ڜ����5����h�$�������p�rVs�X+ `O�9��+]�0fx��O�>��;*�3<a{l[��&�;�׬�q�JI��|O�>vZĪ�Kr�1xS�y�)��1C�Np�����MC�B�峄�2I#��V����&룄>F6J�Cke(��d�a��y�����q��B������*(ci�,�(�'ێ8�H���JkC��`���5y-�ԍ��L�*���&o�1�9֊��yZE��`��C�}k�e0���)�t�A���Y�;v*� � �g� ̖�:ǋL3�4�ڬ�����OJ+��U�0�a�]a�aw�����{���{��r��nF��vD�TD14���E���.�7�>�\D���j���T�t����c��6���?L�*��SićXs3x��E�T)K�1X�����+D�܌����63�:Q������|qP+��,Z<� s[����5:����>-F��,0� 4]�	�UO�wG��\��n P�� ]������QR' ����5�\���8	�Xt�t:�۔��/duثS #��,�o{k���%u�(ǚ'����➁�N�VO�����$8��%�� �~l=h�eXȻ�X-��!Vy-��Js����!Z���Wn�H|';��s���tz�0�*薊��@�X���b���e�f���1Y�q�X �𭸴衮W��U�LU*0�дv��K��|�X�Z�-S�5�>�]Us>�1�LQ�Aw��]�|�K#g4�ɹu\�Fĥh�z����4�F�!K-#�BE\�7�������ޯn)W���$?�����B�Ӄ��^���H�q2������ `H~�4�s�}��b�<���%�W��b�������u���`�Q�+G��q���˜o��|�l����6����c�x�> y��G|3]M!�\�??=*�z�M)�c��M%�������"SB��f�VK��ŝ%c$=n��Y����<<�^N�:�聵iDI����A�r,������pfz�W���[�X��g� ޏ�zG����.�(�{�'���&��9T�>4��汑��v�.�,8�`>L�t��?}k`7�	]�=�q���Ά*�rx;��4�cz8�o
63��$daI��H���_`��A�X�%�d�V��S�'<Yb��=�t�=�L����� ��y�ހ�E��9s�
���zO�0h%�[����]��k�ֻ`NR�$� r_Pw�eO��m�s��T��)��e��s�<�G:ߞ�6��$��*Bwr���g9�C]�.q�b@}�2���VY0%���BpDjz��2�`y�O��6-0�Ų-_�?YX7^u;G3u�x�Y�����1��ix�~(5��34��L)�J�һ������1GR�z"��r2�"�R�7�c3���3@>��h�PJæ�q0iL�m�y5��W��⟜3L�5URD�eZ@��`��yZ�'�E�88�N���]f|��%��A���4�8j���I��t�M٢�&ʀ�|�=#�'6;�=� ��������~����%D�W*ʣ�- @���h]��Vv9���K�t8�_\{i�RV�8�w�;>����E�]�v����ᤢ��ލa��ﻎ/��Z��wv��s��[.��,�$212Cۇʧ��$ dӻ�"�����%CX�6cڴ:��^����z�n���Ym�g1h# M����>qsa5PN����98B!܊���]@��S�Lã�B���՚r�_�2���U���]�ٝ����u�e��#���á�)3C�R+����O�����7�E���Яe��ʌHb�)���~��{� ��9���'��L�b�.�8�2�b1dk��iQ�񥣟[���3��4��N����
,��������&z�]a]����y�`gz��=��3���Ci�_���&�8y�	?G	�*���@������]j�~ܴ��s��
+�����\%�4�����>�L��`�.3kG��#��,i@�����#�ܿ�n��o�%�N7|H�3�Tݗv��:hpr�,����o�}'���
<�4�>@!�ƻ���#�Ԃ���|�V]�����e2���	��^ttf�<�0�c�,�!ԙT� ,�VA�^��+������#� `ug���N�F��RSh�4��)�Q��8"-낻�`�����gD��B��k�\?��M=���
-t�P�R:��K]�ob=B�["��?y�*D���kt3�R��`ve�
�H�`��WO�2i�8�&-���q�9��]�j�S�a�ͧN�6$D�z\ �Ο�q��	,�:!��m�>U�gC�=Z��͢ǃ��F��ߒmR�3�m{uAZ���vuE20�L@j�b�T�qd��3�����o���s)VG�����ّ�z�$��kS�ɤ+`��Z3C��c�u*�Q� !z�ra:���0��%E1�;�>��)�]��~pC���:	��4�ʷ�Aݭ��oz,f�p0@�i�-%+7[/�uJ[���@!����Pg�2!K-�}S_dי��=��:�+��Q���1�0����#+Y�H��c��'���^I�������1�ז��hgŹ��Fj܄��.DC�/���7����|�6d�RWӈ�.�b�=����KǓz?be��~W�3�S$0���[(~�s��#��͔b6�IT�/<�D�m��_��6'`
�mSCC�]��x]�A�z�ȭ`��F�8���
l�����U��Bb�F�yq��U���CgϘq��m�眧������P3�j����G��g��w��;*<,�3$5o���W������mj��F^�d1<��Ɂ����z�O��,�80����)�n	%F�{M�|��gv7�U�@A;��(3�F�"�R�18���|�2yii,�/�U��}ە�̯����}a]��q�U�_)�^_�3�{��dp�5�'�"C�T8a��`D#��55E� JZ����E��;���7��@���}%c�au�~���`ZU�@�"�M(,s>��0��bT�3��4!��#������Ï�[�;��'��l�!�7��e��#
;�!C���ZBcJ���]N�@y��6mCp���ľ����\�Q�~�IC1asӈ����bi��W��
k�3�4�m[4I��!��O羫֋Y�� ]>��i�Z����n���3�_/�5p�"/Е*$�\�?Q��|~VX.I�p��"��dE�
gk-��NT�\�ך�僭"��8�IS�M�ق!
:�9Zd�'��J��%f_�aM��<�ͧ�.,G�S)���X�gWj����Sً�%\7�,�Ia��'��\����@��}���9�of���z0�U@�m��dCu�[FF?�=�8@٪���%��LK��4:�]�d-�*���ʚ-@�R�
~)I�oك��1!�q^��H�rʴ2	U� n-�43ϫܜe��}���qѻ���L&�����(;��tL3�_/N�.f�P,�/��h&��c��߁���X���X�l%�����ܭ"p��˄�$���]��-˵M=ٿY��P�	hK�;G" 7|>>Z���FHM6,J�U����Ws���T���x����k���:zj���6x�R��'0o�0��d=��+����TG׸X�od{�y�_j��y�L V/��/s�xEo��i��s;���!׮��~򼑃)���%�u
��h��Î�3��@d���ܹ�}��'�Oţ���D�w�pC�!#DaH�s�'�`�]��4�5�y �⬊�D�,�K�0��\;
Q��lYo����I���Y(��!�0���r2�+����m?��,��xԙ��Q����H��`���teA����l��	��u�)�Ϻ�Y쏑�F���x�&����zW�L�.X7&���м|&=~tYҰ�70�Q��·G�	#��gRr nԗ���j��B�2汔��N�C+"^���1��t�����f4j{�A����`����Ww��5�����Wh���B����(*��"D���������b3���Q�$qƇ<7"�g_g/&F<&�~a�ܗz��ڜ�M���"���ӋS���(��Ο�4�@>�����?��5NƤ�5�����_�?��^��ق��%*��y �_t`�K$ ��:�#f�ռw��{KF�#|#/��J�(��(x��Y>gA��9iE�Z������W���ph���l�����6#/j��3�H�(�����ue���&�0��s=FXGT�����/g�	
d\''�iVV)s�ݧx��3��zY���lqF��O�h�Z�[�P��1K{�G`Gu+�ߣ 版������52n�*$�Ȑ�i֏n�1����I��B�f�?pI � �Ջq��c6����$��	�cz�~�P&�b~P��+�F�j��څ��f��Mzt_�t�Jޅ6�҃�����l�0N���j�o�uc�Ё<C����I�͟��ޏ纇	TNm�8\�h��vO�zRI�׭�`<].����BZ�6�� ��z�:ڑUڑ4����Ł?�gF�	� 0k�_aF���A_�HQَ7�l���wL�U���΅�\Eӕ#^�v0�s?,U�o2���)�CHFo(ݱ"�hԷz�
��zp��춦9nfGF�8xK֓~H<�cT���9#�i3	�М*u8s	�O��@�i��LȚ��d��RB)>�.�W#CS8hS��#���`p�҄[�Ɯ:�/�������6�T�]����yo�³������ ��W9�z	�|"(��a��!���V���j[[M:�����{��4��u��'��y��P,av~���� \ww��6�K��d�q�s�sr#\�������h��4$L�i!ws�7?B��I�j�^��9�3�9K���8��fplv�*��;TV�hZt�v�L����W�	��e%��J��8����6GLïF���}dr�#۾��F	Ϫ��kf�S��G`?��|9��PM#''."v��s��E�f}/�QyK�����Q�y���z�%H�48P��I��3�e��&^�z:ϸ��|}�(u��L���<��¦x���x��o���m_���;m-��E�7<�|S��}�
�2�V���q�������'�O�Sh��%C&}N٠D�����G�g��Q��1�p���Ё�?�M3��-�����P��7k�Jt7��PC�w�Œ�N�9DFڦ�,!�J0�hi�|�YN�5�X�}�*6��N>�[_��U�ض8�ۺ�;݊�P=�QǪ�2�:6k�\/���6�hAk��!�q;�ѰL�ڣ/G�P�� V/��r��}�cc�?�<<�'d�s�Ǥ�ܴd���K��R�8Xy�yB��=-_]U����~���]��b��8ž6w�@���Mu�1�����mxzFw2��+��^K:�o�
#�F�6dQa�PRmE�~N�ir9�Uw)eO��~[^����ѳ���ٕ����= %}a��?� �P��Zl$Wn� �B���v��쳪��x5G�S�"O���|�i�D��b��ة�X�*Wz��5�a���)ϸ��$A�E��[�����������kǵ�K���&@�D+f�^V��6r��n"�r����z��k��G[�M;��T V����)�.���p*�%uO�c��3(�-�;�k"�8y����P?{>��^�ⵎ8��]_S2i�`7�rn�,�^!����.�����d�Fr�b��ig�Ϳ L9��N�/����9$#:^��Q�͔���glS2l��⇡�婮�M�^N!��j�I�x:K#N�9\i�S�bqUh�n�?�����J%���h�fViyq��]J1;�'i�c��N��5���	t�u�(��ߪ'�:A����Ve�~��+��u�5��3��k�oՍ<Bz�+t�QC<�bfͭ
�E�����������]��rT�v#!�c�Þ�-[ؘ�U6nٮ4����`����*�����P��i�,��è�F⠔�I'��8��8y�v�;��P�5�C�#�u�����޿�y�GrK�/��b�����`m��e[����<�j�(8�59~s�RZ�ȧ��J/��&u���q����3) ���Նr#�ڔ����K�#����g��̩?����в�	�C��R�����щu{"8��Ob��0�N���j���F�/ɸ�P4C睸�ӧ�J9��R�]1��j�8}y��k�K>K����&�B�/`n���V�A�;O���M����8K�j��<���ϙ�mH�d���w�������&m[EJ�O�-OE�~>����uT�du�W\��U� X�N��c4���pi�L^��@�9�2��$�H[8,4<t���*d��h��!��d�?�%G����x���@1��#�Hc6	oJ��X�JO8��WFK!}c��72�(@`� j�n�t6O���.�`���"R�J�y		#k�і�1;���3O-�mʋ��������8�k=�\'��Y���k¸�Y��Ӎ�����������K�mn���;���g�b`?�8��w6Fn�NI���|ƪ�Q�'��Ϛ�jM�M�Z������6�� B��4�c���~?Q����ǌe"\D%���e�J��5���~� x�ƃL00�6=W��ݜn��\��}�w/G]DF��eC��9صn�W0"βcaG0JuمQ���T��-6T����{�TǕ=�f�A\b&e�w~q���8�a�	&~d埂� .M�w5\�E\�#�K���3��{�
��\~[�D�ׇDT�_l�q������H,H�k��"����W쨲���ŷ|M�v�a�ߩ|�Uy�W=c��n���4�xb�q,����e�=�?Z��rIb;L��ɜT�#��$r��<@�@摰���43��
�V�i  ��i�ig�[I��w�1�k�[����K,c=����;��,^� ���6��~z�2���S� zM�������yݦŏ���̖N'�D��Ε��WV��a?����w2��wk���Sf��HD���7Va��D�^,�2K����8�(�v_0�ct�:�e�ؾ� ����P��9JR��ţ�? ��	�=	h
bC�̡UD)!t)r>C��zOҞW�j�L`�G���;�H�
 ��g/ql:�Y��t�����X��X�6!0QV`'��1�����pt����9������ҏ���L��/y�;�����IACT
������� Y�v��j�|�2F�c!_S����a,��Ǆ�y�oz����D�ń/2�rU��O
	�����P`��(���>8@o9� @���ֺt;�����H�=
c���a���� g�`A������
����}���y���ܕʹ��˪0��t:�����<R<u�
�8���ym�Ā��Q����hx�+Q#��+\}�!O��RV���[2�uN���t��K�}'�i^����˾ɴ�;@�5_�k _�D��6z�L�������W�Dk%�
 Wg�[���r���9��}���ȲP3n�j��D����M �g�Í��D������I�l��"q	�h_cP�A��TE;�����^٥YR@��\�{�O���~'�va�R#Ц��*<�oV4kޮ��P`9�j.B��i}޿\��F�v����xΣ$���T	��kOf��cD� 9��fI�X�.gv�����3;����>�$�3�<8})Ȋ��K��5�$M��O�Q��F�՚�)����΄xq��U��"�F���XO	�e%;��Q��s|b]t������Ivm�b~�P��d]B���J��jb�6Ƚv��<���F(�q�d+�M��z-4���aQ�P$'V��n
`D)�.k�w|��hLe���Ŕ`lt�Pܧ{ٔB���`��^=�_ ��1�{��mꯣ}��xR��!#�E7Y�~�ށg�vh�ώ��9�������x��%{��T]��.��f�g�\��t�`�Qr��ߕ�J�niOP�hN<���V2润O{R�*�$��dĨ�a}��4��)��,Ny��ʒ��hI9�[J�(���M_�����1e~}����Qo�te�Ȁ7�R܂�ٌ!�PSЉ�x	uHu�/�����j��R�gy�r* ���*Z_���A�!�����_�%�����
k�]=��%����n��T
�p�ۤ-P�P��L3x�Wi��52��=tL�Β�������0_ǡ��;�q�ڐ�;x�ssYO�������B�����A�0^:�΄wJ���(���P O<�확��]PBL6`@���3���Tn<�`�N��o��J@��e�G� �����Q�=\�m=k3:��0���p�}e��3��������!�1���!�f�]ɭvf�+�w��qT�ؑ6f�H5�MU�A;�GJS���.~W�H�A�7ds��~�l��f[�\�����؊�q3	���ytα�M��Øz��;�7���`� ��č�W��k����X��m{��d&���i+�`n���f~����'ȷ�'�je�{1�&�P$�����'��70sc�����{�gݗP�ŷ3�m 6������*9���tZ[�,��@�ǌ4Ww�=1r�3��ַ�c?G&1/\���Xcߦej|����$�wM즍ZH�o��.�(���6����7�%��z����~|��"p�k{5��F����.��K�V��AIՁ�#�^p���)*6����E"J����u$��ޘ;�ȭ��<Ų�'(`9�ߑ��i_�7�5����
kn_��\�;Bň�ʤXp{ͦ�`#�O�����O/��:Y����N+Y������F�T���ThhB��u���`ֈW�&�A^M�>���߰?`�A(��������c�Okv�`֩��{�=����01�ϥv��4z�wY�1A����h�Z�!�<�Ag|O��e/���qrH1�0����:�¤�tXa���}�D/$MS5�<KTu 25��)�jSij�����1gE!lb��s�&�B"��T�(xmP���a�iK�+������׵�����3�X�^�oY�M:�#���o"�Jc��9 {@?��X��A��>Ix"�~��y�?�7�6���3 ?�����@9��
P��y8Lp#8���\P�s�,B.�0��V�(�!���5�[��1$�d���/Ѱ��k�-d�V��x	��@�5����Q�Z-������`J&D["E�k#f%��+�����D���0�2�P~;�E»�9	��>Ww�a��L��U�C7��wmB_�
�Z�b����$�8 L�����|tQ���Vv-s�۟�����I��) %H6���N�=���k��}@f���ʼ}cLz^�?juz�j�~B�*՗������wB�yK���I�3�=���5�9��H�d'���	��K�5 y�M&�;W��站��4����+�?�G�ju�'+in�ac�F)�� 2h�'��*c��G�3��h��3��[�c&}�P0`��̡aǮ�绚��>���8��2]JQ�ؓ^o�� i�Ϥw��8����p&��ߚ�ǀqj$K��1�0,DI�E�s��5"T%�InF�M*��)�2w��bͽAȉz����"�r�{����l�؁l+��2�+�w����������7~0lD M|o��&��I2����N�7��E$�K@z�ˬ��	b��[�K�a��ǅ�>LC�;�
ҁ6ݨ'mi8�e�i`�S�ψn'�k��S"� ��A��q��1�wnۭ��#s�ώ忩��.��U:yِԔT�cK���ic� >��b΋%�ϥ�Wr��!�jp�����c#;~�R�ň�ߐe��s�����;h���`!}���8�t,��G��8����8q��Kf
�GB�����c5�7^���AuK����Ab�-cG�\�`�E)��9���ᜯ!��f�����Xa�gC�<����{{�)z$Ӆ3���F�&A�e�?��(��K��0!�=���o�7a��l$ 9'6�mM����ω���&2��_��$h�"H^��<�vVt�J<��K�񸏝Q�i
�E��c*�#ňv�9�� �>��1utg��i"[�p����G��y���1ީ>�[a@��%Y���=[y��FvL�A�������W�}Ӈ��7���I��vuiz�$K�0K���H1V%?m�JE��� �F�����t��~��q�{?����g�8b��Zm�z�;�S��N�C7�;��-��
� ��j��V��Sݍ����g4�)�Ls���L�*/[[2s�������}��ۮ��'ڮ�a�خ7�e���3���|v�
����|�PO�\G��dR+|P G �m[<=r�2�UZ�����R�����F�DY���a�<	p���cY��q�β�n���r���q�N�Oe�ƺ�I�̠�����,�2emSӸ�2Q�N��b��>�al[F`��5��i/^G������P�4��O��U��Z#Ip,��P�D�7C��S���n��3��?a��Gà���m�
��y�:�����?)#�D�ѣ�):���j��/�'T�Yo�Z4�2a�<n)x�j��õ9�;�y����aw+��Fc?�G�^kUh#S�&0�fF��:���I����wCt �wb��5q��f����� bkOu�!MGN��/��Q@C�(�k�Kn�`�����Z�r/��1���4�)�}��o���6\�=�ծ\.�F�:�SAv>������[����Z��0�v"H[�{�Y�M��E}���,5�MǓ�h
��P��Eɤh'\�U�L+����ڄR�8����t3�'%|X��2>՛�������_����2��x�^t������?���B`PP2@�;O\���҈;!�mzs1��-�Eb�	�5Ml8?�?^i��^ذ���f���5���-q��������0�Z�I�����Ncp����e�bo5g�;�4�q���n�Q���NNS�̀?�k.��⛹�$�aj�P��j�١���n����<<nw�z(��38�VU��;��*u��R�47n�{�� Qu,XU�ua �h�4�8%܀�c���ֆ��x���>}A��֒]�
�>|b;
	,����8T���ҟ�	2w�|P��%&�/A���z�7��m!X�T��3*���� ��	c
)�Νs
G~nd�2�fdZRIZ��I�uh�j&ɵr��.��+���Z*�ȫ� �u�{���&{T�'zR�>�K�y+�C,�	����V6��5����UL������>�����,N� _�� �Rp��[�A4��e7C��Q�J�o�A�;.��ڲ��~I�p�C?9��Sy�)��ţ�|�-9���؜�'W {>�-�g�ÌAɉ�f��>lex&��*n�H��j�7Ҽs`]����*}���Zs�^L� ��>�A�0��{�;�C�qƎe�jW����{"��$(����v�m��Mv�Q�>I�`�jF�$�MNEg����
sZq��,��-;J}X���*��3�
��b%-G�ZG�~xg�f"��������}���K����6m�c��E��7���I15�"n�-�G��{�}�,����V2 �Y��C�/\��0nU��^�)RD�T�ωB����I)�qR�`Q���̵
j�DJ�����Ӣ{�ס���#1.�4ғÀ>�"�Q�ԉ��� �� 9��맱e3�=4\���8�:ZVQ'���!	�{�E-!�i�G٭"�'��Q�w���Z����g)\�w�+�xzc[�aE��x��I�	���8 �"���_�l��Z,|5�!���oj�h\� Q�J|T��x��s��PR���}h@Җ`\�{�9�Ѐ�� 	w]\Ú�MW|y���k"�j��r�^8���e�"}�������%�ĂN}I���}�.bcx��+�2�=�\�+<��cM��Q�v4X�ǘ4J�e�LV��&�/�������cM���a�!ӣ�6�="M���l,Z��i�R+�3��^fH�}�Z�MPa�ʌ ���eB&-G�i���9�Y9��..�L��`���޹��!{���i� �@�KqO(�^+:xB����]ֺ�z�F8�\Cj���x�g�d�f�qB�h����ץ �J��9��A����v�9ؑ��O#{�T-U��\x��P�?��#n�Z~WbX�U�˷s��k��z'�%�pИ��e`�:��G��Q�d�y���|t�V4~��$es�q��ʭ�FG��MR�P�a؜�+��e-"Ea�=&�k��b��za�R����2R ^����լG%f�f�ݺ�? ��$<��C}���vU��N����<_�:(>����������6����/O�4g3��j��Te��=WO��e��&�����妀�>��q�ek����|�݈� ����RJ�I�>��F��_�g�>}�x6�\ߪg�9@�����t>� h*T;t�T�l��h�Ǿ�j.�حmU�"�Ynb΢���$wQ��3�@�a�PA�̽��.h`t'~Ya��2�=*�+�}�� =�`����GϥT/~�ƀ=�/D��~|9�q*����R�ДЈlJ�G}��`qa�������tBHU�����ݥFW��{��u��lȚorG:�<�{���(ĢM��s���o�#�儰�ʬ�A�kg���y������$�Ϊd>OS��3���x��c{ͥ;}P�gP��obp����0�W�@QRT���y�t̗	c�g&u�������(�iM�R����S$W���֝׀{��Z�$��� V�E�7�����%JJ~Q����I��wj}f�.�0�.�8z�a˳���7v@e -7��?�d'�]������'���&���ʉ�@������,��{g2_QG�P[���x)]��wؿ�J7�҅66��r2�WY��+0���l���+àl_YQ�J~eV��4ث�U�e;p|��qy�h�u�e�6�w�P���1���N�ĈC܎���TM�������p��_��I_n�8?��CI�3�>P\�&O>��
�c*S���#���<�J��L'�k����3�J�oh]�(��R��J9а���zt˖4�Yܡ �<3�l�-@��
��m�}�d�=I�������g�Y���a}f�=�Lv-#7���hK����x-�ßS~iG7�4tKL�������hҦ�-%q�Lp/ ą��(r�m�dJ��g��!L[�h��<ӆ�R��\�J/�U��X�OA�}�M���̣o���h?Q��Ё"kR����3��0 R�iId\$�j�񊒸��RqM*�|LYf�a,/��6�z�@��*�M��"���Z:k�������
u�,�ux马�8�Ǵ���b���5�v�ʬj�N�N��6_B�E~C��I���L��(.~� �?�@�Z��c�[�:���7H���`{�#���Af��e����Kr�����.81��^��S�5��`q2l�9�W��%b�s=�ͥLa���kݩ�2&�ܞ��IR�;��n�T�������ȴؑ5�&�� &[��5����l5�U�Db��_㛥�")m���s���<{؁s�
&�Z�>e�R��MQ#lìLIѧ� bo���|�>��+�X�������t��|��Y�H��X���qY��;��LRE���́,,$�/x+��K�A�9��@�5�.�E���h�r�|4�}��C���l�87��=D���Vj�@MZ1U���(e���c��i��+��I#^d��O�zU`�u���S�"`!�)==�b�V�D]��j����1��O�$���~�i�%�׫U��6�#q��1ܝ�d��b^�&G��z�+�vy+����ԯ��)&^�%LU��Nh�4�[��iK�b�2� ����W-K����[ p
c�컍�� �Ʒ9� 'L��d6c��ٸ�}� �0+����P7}�k';�g{�n^h,���5Z�i��ԓg�M%�����Ώ>���p��n�%ul�/�C�~�ɋ ;t^�l���wC���s	�12�Di=0�5�^��k���d׋\����;����Uhb�J�~Իه�ƈR� b4�%S�t5�oӮ�!O��E�z�n ����]:y�)��TFr�������&{JЩ9]�����:a9����ц.F|F��ߓ1�]�L�T�0�J�!nЋ$�_���dy���r1�
�
hM:��Yɞ�̸@ڞ:����Á�{���!�,��a���o�x�!yS�,����w/\u]�Q5�'NnG���4��aۅ��gx�6�F;>����	��d��⠷�����8?�������V�o	���ɥF�?��L���������Yxoy�I����F"с`�F��O�8z��(>ء/�O�;	<��n��?�`��t�#��Ó�.��$Yp׸�ӌ��JeZ,���6�	��H���tW�<B�}�?�����0�� �˄��.;M�[�7YF��OƓ�L�W,`�m�V�,*���J��;�d��K�$0)�6d<[��e�b�a�ڃ8���Ѱ�}g�R>�}�tf�SA/Nv�SԔ9��;Iͬ�p��P��}J<&�N��O�wUF�l���]?0���`쳒D����n����� �M�1��gؘl���֩��[�(��q�&BV�yFŝDa���/��B���B��7���z�����ǁP55x`�;������l�`�{O/�^⽒s��x��P��`��B`6Mߍ(�'ɇ��! �)��C3+�	��2x�
^ңM�SD� l2�����C��t���9n� uK�ɿ*1��]�bN�w��coP���)�&=��jac|��6�.���_��m2�3W������|���&����B������d���`>w*δ�?zvo�������n
t�XI����}����[�0*,�Op^�Ѓ�p�n컚J���#Z�����=�;��ӂe��JGEm'��K��C�f��ƎY�"R�1�Ș��O��Ư.O�+��%\���P�;F��[���\#�����Jk�lB��<<6���~�,� ,_�����g5MM�r��Q"΀Xi�MF*�k!I�|���,�@_����RIm��}�<ۑi�L�ord�*���a҉��� g��C�$L�=��0��1�H��^�i��=#N���Bt澛���*��w�DT����b��-�y){��Z�={�$�GA����*_ܾT����Й�Ÿ�4�)��&�bq��Ay�9,bwR��Zm��R������\./J&�$����K�Hj���Z��z����ɋ���:U3te9PKs��n�𳓜ܡ���T��T�g�.P�"E�ͥx}��m�M�~�lC��%�k/�M�/zk�Io%-wr'q|��(9��B|�c��A���Y�=c�/�j�����;�".�u��ʾ�ed}��%5��
/㴧�X9��Y��`��Өуs?E���Z�-��Zhfa�3���s�+�f�$�{��^�����'���X8��R)�3����7��Rәf�f�P�>��qF֛��+��-�	yd��1��]�jn�ls�w��ļ�����	�b��Y�P���8��0����-��+�S�~�������6"�\&^�	�$���7Ş>�������勬 ��^�Q[��A�9<�B��������&��;�O��r��l�T�nuU���9L�w�&��̮���)Il'9�[�Bō�q��}��yn���װ�|D�>$`�ag(S?�8���j3���l�0�P���Y����|����e!M���"C��\��;0g)�����zD|i�	��B�cd�>FRmK� _�~�e�I����a3�{5� [dB��bw� >:˘�&2����������ԪCQ�(�x���b����̹��b��A��Hv�̜�&���m7��S�����M^{�d�/+m�Vg�\� �{��el�]���$�4w3b���[9��=�Mq �l��4��u<���΅���ۓn�3���-�*�ۮ uWɠ�K�M�_k���b �C�\��X�lYVCT\��l���w�*��
��1�tK�GJ2�b�G��SN��oZ�v��d=��oT����>A�rg?E�S���cư>�ck1��:l�:���.e�Jej����j�����q��Վ"�dјVgĳ1k��������L���%|�o��A�cOh�c����g�J�Ј�A������?s1�D^��^Axw!�y��~��_�vԋaE�	c��x%#�`�;E���bVU1V[�g;"ŝHl�X!���(���i��]<t��8��#W�L�suT��V(q�U�
eZT�AC+��J�|�eZ�".\oػ�>y�e�2���3�ֵ����O���#J�?w��X�.�׺樛��֞I ��2\OX�Y�~��dѻ����gP�=�e�3<**o��0z��aj�-g�eY����T<[;�� j�m�_v宍x�ӲjX�~�������51_����X��
���8��,�"��~|���`����Y� q���5PӪd6���j�I�n�(
j�ԜN���Lp���\������B��R�Y3�}���K�[��<~��5�~2d��,��t��R���f���'��ٛ.O��ՙ=fzo�_'Y�mbMo��Tǘ�к*.)�+���kDr�pG�[d����u4-Gc�c����<�"<sB4F4��̣��X�]���¯���{g����Rѳ�\��Ŗz�>��S<O�%у�B4�I��iB�y[���fN���|/Ӂ�I'xP�Q:b� �_A��e�_�H�o?��F�W����ZG������~�i�c���'���dqk�����#EY#�+��@��|��A�k�ƀ��鷜��C:�>���'���[�R��<y]�P��wt�S�cpx���-2���zۀ�ŕ��
8�D����2�-��ҿ':jz���2E��X��nAx���ɓt�c3��O�$�����))�� H;Tz��&s*�׺�k�>��ѿ?mE�K����U9�YB�C������Vة۟�W��! h��Y��T��憥a�e�]ԔP���}��� {!��T�i�ÿ;�Ԍ�D�r�ّ�S�S�����J�1R"��,��Y��[��6=�w`���	8�?���<��AAƽ> C/�@7��e9o��,���C�~�W�;bH\�x�+�	f��='��j�d��� &ưeO�]S��=ao�\i��m�S���#����;Џ��9ȩ����F�Dڢ)+:��S�F���Z���WfTQ�hȷåi��:U�l��_�;�󏳤v;���E�rn�y��U����Q^F$�k��9B�?�M5��c�VPbn=>�B-_�z$�d�����4�+j}'7�o�כ�.��F>�sz���T»Qi�\���ƊTX�sl�C�%y��x�4�N�/'�wEP��@r81�2$>��[÷Z]�?{ �T��}�h�PC�"���}I��_|ĻK��*�Y��$Ϧ4<Cqۦ4����$i_�I�m���sjO���^X�車�9db�.��֖O��.�w^��hx�G�M���`_���4D�c������,id`�1���n ,��yJs�G1�YXji�[�o�����m�����3~�U��E���p`�uGk t���Ά���r��^t�-�Yi��@O7�Gd2�68�n�����(�m}4��n��ջ2*l��k����l
���1�qf��I2+����S��`]c�F�.[�7\���[����`ě婝�]�]cm��Gҁ_�D����&0Q����� Z�t�?������*��z��� }��\#�%�?C��+���(�6�0%q�KK�- w�+rN
f�S��q-�YF;3�ۑ��&@mbВ�ar�|��U���^<�:.k06���밹\i[���� s�[�M�a���}zK�L�1�	�.��-�Qgdmu����t�q�<%��~�9��DH"�4�?���-�אS~���PD��x�"*�0�J���&yT?�Y^�q�ߔ/����g$�v$��V	��:���3�[����ll�ă�i	�7�y��C׿3�SL9nRr�
���d5�WZN�[�A]�0(#9���1�y]�&��ѵUll'yi���}b����A�L[
�
=A��U�_����^¹W��\�hj��f[@B,�3�␏Xˉ��{�� *�.0��?�d8�����Pيviu��æAk��@N8�ϠQ
�@Iuj9#��F@�QE;���H\���o�tǩ��<��>vx�(��6Y�Ld�o��q���c�)K39	cv;bWz����O��>��*�T=g��I%� ����u�����x`�SL�Y�/�.,�|g�ũ~ q2FM�\��W�"�{�S�%�
5
/�IW���qs�p��r$ 2�cNy�ر� ��u�T�d�|��`C�{��DE)��X?���SQ��k������7����"��D��ÿ�IҥCxy�C�L�����/� n�*o���,�1�eᶇ�#�-ʲd(<`m\E	G���!#��y,	H��R2`�$.��B"j��%1������(�Q��\k���$�j���_�ޤ�O�.�àƦ�~��)�e��[8L�D��f&׶�������?�5��1m�7*�#����K���W�KE��y��cTUʿ�P6^��Ư������
;��t�I
w�m8�)�� ���:�֪�P�\��8�fK>L��^fx�a	Aeс�G�_�ȥ���X�'@?-p��6<C'5Oz��+��Y���<����w-�y�ߣ�"m/aiVZH㼁�Ud"F���5�2-crnK#��S��>E�������"�^�w�>ƕ>�p5��n�h����{�x7!�f���s9�V=��ǅai�7��L��Է.�Y��OD!N��;�lL�/+�R;_RY$�5������\�TQ�;2d%��Q�(�r�>�a��2�O�Qf5=�u�^�tG�h�VO���b���Q
����ݏ!P���%�;zp�Ðo��~�ɕ���mɀ��'̄� Ѱ�ޝq�;�-�  ���B_~�-��\���6	���b%&ny�me��h�n�\��������� ��΃�`?X_��p7c$m	��C��˞�b����y��I;��<F��Oi�!�. ��*/F�ibLc�q����H���c:�}����"N�m�Tƀu��r>���v�ԝj�O�/@l|I& �t|J̳�%y/Ts��H�?�R��-�1��e
_����s"��$���RP�S4���m�gY�{Z%£.��q��7-�ph�~�R~�3���c���uK9=����� �m��a��
, >�"��W������Y2�"YJ�3��^���r�+�e����>�+�f�*�bd���m��)X6 /�0�l�$G��˚���5�&��*@]�~&�@6Ⱦ����3r���K.�<�(����f�mڊc�s��GNᬇ�]`�n#�D0n���3�A��%Ts H�]����{_�ш�́�:1��Lٹ�/��ci�c��Z��(<<��V^���`£s���Ҳ�`Յ�
N����[�i�=U�� G�3ݤ-����2�#\x�y&2��D�q4H������c��$(Xƒ�S�αF�r���yZ:�~�-P`%"����v*�\�rS`Q
�@�ح���u��RUY[�<�K�ݾ<�~1�^<��_L��r��"w�N��>ؽ�z~�#��g�Y��}�^}B��Ɯ�RhB�#Ҽ�z���S�S�7X�k�nބj��Ɓ��K�����<Jn���a53v����"���tXX��at��eg������)�l�&��U��6��7���6^�*EavSoQ�I�HRh�{M%ts��l�M^}��K��o����f�=ڦ_y�d�2�ֲ�|(�q�u�۝������A9_��HS�9Q�cg}~77U-�������$��[ מRS��p;�Xz<�Dp� 4R�O)����Y�F�����#��&��n�S}���Z�&Q�Cg%)��T�JKf8�O7�>�l>���@5p|֒˰�
�5��	�-�d%���q�xÀ{5$���S �����`.)��G�v<���YW�̎$�\`�D���B�<�gxF�bO)�u�<�Z�P��3�;oA�i�Y�~Z�$�A'2�s!#p�Z���673��p����Mp�ʋ2]������qu�R�UP@��_�A�����3�l�t�J�I%E����r/M������P��Ml��@�k+:��'���V.��% ,� bG�	�b��X��hr4k�|�e�W�{Z3��]G��֬����&=�9"<Ue���]tv7��կU$틀�d��p�`�Me,83hKoJJ.Q7��E�b�����ގ��29�>�6u���k,{�75 %g>�/�+��~Vq���k����{���
W����vO��^��������D8L�'��6�5f�;���ü�^�9]*�t%=��u���2��Y^r�Z���N,:�?P*��O�ק���L�8Z�Ӏ5�aJ4qH���-S�m� )�B^j��l��H�1��E�a3���o��k���E��r�2�u���_�Z"�7�D���%)�bKs?��˒��`��rT����6R�~�l�t%�?�����g�9�'�XDz�:�`� ���U����x�$�O�v��=�����-�M��a�8[|��sg��U*�v�zUJ��Ħ.�H�����h��͐�!W���=�/r��IE�O'�mp�2�����2�ы����QH�"���� �1ƤϬ5��\��Ś�l�J��j�����딨�hkUX�m>�𲛒��"����h	w!<�x7J�T�x�q�2���}8�Y��#�@���:2.���@�ͱ����3g)�;��C-������Q	���_A=p�}3bla�j=ڊ�\�ݾn�����ӻ��	��d��$�v�gGxFX!�VX�)>�M g��ћ	�hȞA��1�b�^l�M�~Xm�V9ծnpO��~�:��u�wf"ȺW筋�9G@a�ɪ���Ri� G��~mP^L2�J:�_��n2�_��`��I�@�)�
�vznr�!4I�c�l�?�6Xr��F`��%�00;>�$�bŇJ�P��tb7���\�K��,50?�2���f)q��˼�'Q��6�.�.�mJ>L���Yr�!)��#�<(�����ՙ�����lO��a\����.')@`�nr闭��9/z�!��o	�d^�2�4��Q*l�ʅ�7r�Gm��C�$�߬B*��S���P|sU����e��	ɲi�
�����U��:;��u��^a4��\��Mͼk������Y�z��
O�kU�����&	�L��k�ǽ��ͪ�09NX"���&8=��S��1�����\�P���;���B��q�,	�S�����������K b�Q���YUD�k]�;I�&[�P8�74�M�<D��y�����kF�h�b�s��vap
�� U	���*���!䌵�*e��Ƚ�j�xm�U?BT��`�ݥ���� �g�|�SW ����F&#�7I"�PJF��_DI��^�/�l�v.m��i�2�:�����Mn7eΖ���1�Sˈ����NL�˥O)����}��_�����G�KRd�̼�2�Y,G5\�Y|atH6��m$�u^�=%�
��t0�_�`V_�lw����	d��=�PN��+��nde�1��qO �.X���`�Ԗz��@��p�BT���y����K���¡�}ӗ�a���n���|��xA����N��la�s�u5c8P��~�z�Ԇ��������c����+�v�.=�uǯv�p�u���/�nၨV���hoݕE�(�?���{�j�+Jdn �����t��i}���crn|F�[='�b�������K��k���#ᄲ��7�=�u�z�7䫍��z\f@�~d���U֬]��'��N+�<`�-���~��"A<>�܌տT��_�@��nCVN��닏w���O!�^i������g���]ǅ �yt������w�.�&��h<��64��s�v�����C�pg���J&�ۏVIdsD�\)�V3��1B|
݋u�����|��4�!�Ϣ�Ogt���i�k����&!ܱ���B֟>��!biϯ�<�EnLj��tF#bu0Y�9��#F�Y���L��[K{"-�t�#~g�\�����w�����1w��D�~xP���Ȼ в��;�������r��0i��o�1���meX��i��sk�EE0j�]x�Đ3C:P����T$��f��A�hN�55f.����Y|�F��zD N��{�`��a��>is���xDĘ�;�
wV��iZ1�g���Q�(F�xm��t���v5�YdQ���,,��N��=�I��J��j�?�+�_ ef�)˹C��D��Y/�b�d&5P��A%4�3��/�u�d7�Y�� �����(��1�$':��>�,@�I���RG0^NdjAm�1���P�� ri�vD�d\C��^��YB��;�K	��p�	in�-����to�h4���R2.�TL�Mql(���b�d��2$��[��p�$R` �7<^}M5?OS��+��;������\��(�=�}�hB8���~��;�ATR��v������γ� ��d9H�,�%�h8������Z�H����s���9M9�Ɯ����ԧcc��W�R�y�b5�*/:��M�����$*XZj�)�� f��<}�
\��������������Nק�G���������%��ˬ������,͂��t���L�t5�6�lWD+��I��ܰ�v$Yc�V,�|S^�+�69g~���	������jh�	+�M͓A�!�����^�F�?O-�b��?Eg�Fw>:,�0f���`c$�or�ك��,%�mW�մ�}���@6��|������[���zl��z37�a-�ӡ6R�KXL���Q�3׆�A�>SD�]�F���X��A���Y�ނ��S�XJ����|WGb�L�\g(�cd%o�օ��B�cw]z|�� �L��Sڮ �f�}NQ�g��ϝ{�79�$�g�
s�5k�"@ݘB3���^�Kc�s
��sj�:)�:�^�I�n�
����j3�����Lg>�����{�"�݁5�뛼n�������F������`���(��m ;��vdyvœ�[�F$v�=e0�8?��>�!9}D,`z�����Š[/.Z^4�9/)E��2	]mu]j�a܉oa.��쒛����:�V��R'b� S����;��N0��h1S���ǝ���_\���6���NF�q�����j���YȰs��B#�g�p�[��ń@�N;�.l#����_<���13���dD;�~��_$����w�Z�\+�MN����W}��a�����f���D/��>19���� ����)P^l�g�>x��b�\@��Q� �5
�7`�d��%���}ڥ��ye1����y��~��Wlt}�ȓ�?���K�a/������Z��-�.�@���&�6VGc��?�����ʀ���F�9�{�Jx^��(�d�X���Ke$Aץ�{�H�	G�V|/�
x����L�Sm��o:�ȋ}n){���J�)Z8{�]��0s��kn>ɢ澜��z�LX�#�$C��{:���HŹOؾ�;QIQH�["f(5���/�_|b7]��I���Q�O!�I�</�c'X/к�A�o��-\� �"j^�(x�7�n ���D���6���&�WKQ�	�� ���.b/9����{�%��O1�6پl��_B]�Lc�:?wI
�sL���iA�kl�#*�����plA�vz,�g#c�I8� x�f6�����j>.������^�"�fT�k��s:��_Ww��ɥ��Y���U_�)v|�Б� G8%��g���6� N0�ѷ�V~��Hp�^U]��G����m�S���v:�D��A,uX�F��|�����F�?�kC]����9�4�Ѹ����=s�����@o7�p���Mf�e�@*�����^���rI�Q���lbߝ'�=Hhi�$mP�̇0q�BϋÖF�'#���}�o�0wޓN�4b�l�rP�~�p�,9N�؁�`̧��-}�]���LC��/��x���"���sg�"��ԧ.�^��=�:]�_�T=3��L��TIdB��ޗ)\���*v���$?����{3͠������؇�����.@&LMŎu]r����%�����,��|z��&b�Z����NVP��Z˩�GJ�6�G�7���
l:2a��8�UdZ m]�a����,�}-�%���R3q��k[�Yf�Z��R������vg�`�p����ЫM+ٟ��$�?7Hx	>{�Iv�ZuA<2E'�-gѦ�0�X��{������(�dz�c�����������;�PKS1u��'�dE3NsM"��d��J{�!�$�b�"����Jʷ$�(��1;z�Z"g�x;Ϭ�|�7�V/{ixx{�p�'��׏�Pl���v��u�ʠ��#r���q\�4ݏ��dϿb}��c���I��ۉ�#,
�V"�H|B��賢Z��Y%.�b�i跣��Y;��n�b�{�Rʹ�(w�KP��#h�ζZ�9 ���4��WdM�����k��T�g=�z{ɛz� ��47��LIS��]���r�|K�3�#�.E� +�+N���)�Pfb�+|�M?w�ջ�]�n2��M��}�=7������C?����3@�\�D��-?���D���Eiv��,1��2r0���3g�A��qW]�\�#J=�8���#�b#^����8�A� ��_����rh���
`1<�R�B/{�Ȥ��C+�^�#�ftkT���)�v��_Kn2��vΆ�o{1����R��	pxH�ެv��P;Z�w�ߤJ
��g4h��1����p�WxGѿ�����Ts����:4�M�տ�nq�Mk*
P��K.)�X�1J��jdow[�,� F5�ے��s
�"���L9`�C��9G�0��Ҿմ�[-U�Й�n�x�Z�k���}��	�fL6�@���w�͔���ܶ�lo���TR�83F8r��9և�0���T��_��9�Nj�xK��q/nܢ�QVc�hfO���t*�!p�^a��$�͹�Ze��Y@g����]V��>$AIx�͢V+�A��'j�,ɦ<�3눺\0 7IG�h��5��5鄮�����?�1Q�t���+Q���V$I�遁�p��t��� �U�/g+��*�Iz�2�S�K��@1��e��a��y��S>Cp���DZ��P�����ʹ�xg�@t����Ҫ�lHx�1G�m�B����+�Զ���{v��h���	�c0�ٖ�E��+����0-�_�j��h	�B T���O�	�W���,b��r}.[�t.6�GWS^�&���5j� j�-���0��4-��Hugk��ٶ�
�k��~����W�����x\<�����V������<)��^��K���)�8�{4���b�cms�~�%�2k������k*H��	��?��BM� 񔠫�<�&[VG�/xH��C)�}��k�Mr]��ٸ��ʷ�_+�MS�r�U�E�����C�H��7��"ץR�6#LHt0i3%�$#?p	%Kn�.�׉h޵����g�S�������e�>58�?�B�����<��((��B�{j���򟸝p�9ݨ���] �h*��F#�7=�Q
��cr����O�����
��b"SH�@�8�SX�;�#���(�~�	X��-�喦U�W_Չ�uI�X��F3Y�~��$�u��J��7���Zk�����=m�{Y-:��/>
�>F�o�׍�����L��W�a���T���?9�n�TR 孂bA8Uk�?�ek��I0��Dk��k���s�qֲB	c����$T_���������{I�@��!���jKֳ֐2xR��r�}.G�2uL@k��Y+%��гBEr�~�Uy��F -��ŋ�j��{��� }�^���p��}ߩ:ȯs"j���(v����z�=>�Wz�k\V^�������_c�o�b6�q��WU��J�B7q��C2*�ls�~�T9J��m��2�3��f��e�<̚b��T��4{�4�[���/��1Z�U16���ok~@_�]=^�^���eEYd����vp���²V3�X��F�8fS����Cw�����j.���j3��a�k��J����5��S5���8t�m(�
�Q01��_;��9"�5CR�l�{w_��~shJK����ZW��$�g�����'9w0�P[l\���*���o�g��]\��d�f�ƕ>N��L���F'fM+���(�d�敛Z
��Ũ��µi3�R����s�8!��[�CT��c���I#�,��e#ǩԢ4��m����]��X\Du��m3���Ԉ�(��mA@����&f�*w��;�����OT�IH���g�� �,�����B����Z)w������P��4�'����
�z0�%)WD?Q�)�ؗ�ʖ��v/W2�F��W�gԊW7M"S�R7V �`hE��G��U�����yA;V��{U�SЛ��ա�i�D����8�5m>���O���޳���\DTv~N$5�N+���=�Н���/�.�ǬA"�1pO�Ng�sw��J�b�n1�#��NLE�@�w~S��ق3v�]�	�"�_��M�mo�V�c"/1�+���N���PZ�{Υ���*��c�b�?I���Zy�/�K�/	��wreoI��X��)�H�����0�j�ԛU�s%�&�z���՘����I��[�
��G�_	&�Pj��U�+�������u�]����pz놳
�\�o;CU-?�2��q�G���E�}���ݳ��#Vn�}kIP��"91�����7�!]^2v�$&�.�[�u��^~wV�I®�� Vf�G��nޱE�'O	gH(+Ru1�6.<~�W�ݏ���F�?�
����>\ܥ���6Ő��WΛt���jY�,��Dѳp��2�A�ؼ��5`�t��o\���GD-����֜�W���J�6�uvy	�Cx{_P���xB&��'px����_J�H;�'�]��`�S��{�b���d�D2��;I�Qƪ�S���mA�y�)��o�E�>5��9Z��r�������&��xw�pG��~(Xc���2o�& L��y��'1օ���Z��:#�5ƈ�����[bVF��t*����/���ğ��D�����v�:�A	�LI�b]���1ѹ�w�������n´�P�i:��}��-�ܝ���U���Ջ��>B����/���44]��:]�J,QE���<�|V�U�)N�v�<��k�q��a�r�d���e:z�9 �xn��_4�YT�~�pW\�ue [���뒮ïN�{?W%8	�0۠��όv��K�u�T��';Q`9��&"���tId�
��,/��^$��D��=S�̖�4���lL������s���ژ*N�&��x�y��Y��]J�i��G�� ��:�ƒzw6�6��v-"(g	����|�So�wS�t�.�)p'��G��W�M��3�R�@���g�#���*�okX��y�yϘ(�8Q/F0�v��4<ҙU��VA�f#З�ezf��eu!�P"�iI�:�,E�@5�1�OC5�['�.����Q_Ad�J���~Bb�6��CG��+8[�1��֮~���Z����絯l��c�񜤫c��o���B	��B��s��rݕ.�d���|�,���e���T��:]W�"n����VtK���P��Ǻ7�i�Z����Oo*'Tau�TXT�!��t?:`W��?H^�����vs.=���QT���B�JR4O���x����K�d� _b�=(\z��Z�^�@r���>�#�f�%a��עe���?QItl�&���as*�8B������G���++�"�[7��/,��ܘ1/��`w�^���?�WG�q%�@���Sʶ�u�QE����y���:�=��!$!�k�鉐��6Mr��L|�C��`���稯��d�Rka�Z�|��>|�y�v��^hyBP�huf���x���,<�xr�K#���F�H�/�?F���*a^A5eN��٪�NI~5I�]��k��+g�AF�e��3}=_XB�W�O�Js�{�WG��3vq8�0�։�;8m�v��hd�ߢ�B�0�V#��a�^��ߢ`
7�E,.�^��ua�L�����)*�?�VKp\%��t���ݫ�����b�}�'�.kYʬ&�$6'O�i�i7p�H���e�G���IM�D\D-�?2����{&���f��ⴥ�4@�{$&	/X�����:_Z���@�o"֖�#<���Q�<�
��K��q�3}��H�%џQ\�����o��o�B�B!B�������rEׇ�����Ӿ� �H��J�����Q�
�ݏ�2�h�ײo��nX�g,Q5���y6���J��!����4骪z�\u
������nb8%0�:}X�)$��.������5��
�Sԫ����Ig�'����gz��-�I�R^p�p�����mR5W�1��qwO��ە��֯F���ܠ�m^0})�e�,<��	��C�lyo,�����T�Cq����9����	�!x�Õ���f���5Aop�.��~��]e�c7MW���/������GPO���ê}�R�Z������=�@h�fh��\��e���u��e�|G;��/{�TCk;qw��V��������mz�wb�qSfZ0t������o���(��­$�=��
����C��g�Ð���փ��T��Z%8��*�$�I�dDp����E)��G�M��_�o���f��o�8+�z����_�	�:s��{�:ӇW��zQ��%İ;�B
5���	f������ɼ��p�cF]�kM������x���H�C'~����4�c����fm����{�����O���&�lg�	���;M�T�� �Q�,/ݠ��~�O�a���Wi���3�BV�P3����M�����ÈR����:�6�3x����_�n@���{y5���ȓ��nv�NƽR�q]��Ϋt�UI���ʲ�4�sh��
�'E�s��t��j���`V,T��C���BZ����G>=�93�Ts��(�W�=�\�]��֩m�[�r:��M�:-�]�ψo��!�J k�`�S�������|�"�d���e�[��k���V�,Q�0lv�,�@��[~H+;�&�s�1�q���,�,_�ȗxO�<�V���p�la�tN�$h�'��4aa�� �B���CC�͊����aX!��?9�:Y���t�� Te���dAZ���IS1i0�I�]$Կ��ɞ�w~,��E�lt�`]E)�:{��h�HF���W^��A�� �ܯ�A"�R$/T�-K��ٔ8��It������Jê}�6� /ҪM=������'2n�s3�5�R�J�QI�\rwԌ1�!�(�2�W���J)
)2$���Aj�[�fG7��ڒ���9iewt^'�2��0�|{h��(s�P9xh�����V��5tQ�,X��=N)逝N���.��3сL�����,5Ʈv���Gl���mał�������$@���"TR������A6�?U�^��H8@�Ry3@���yd�k��9���ϊ)�F|�4�)�cǿUܴ��l��� �݌='hD���Δ��ĝvtnkBi�JZ�l��d��,��H<A���Q&��p#��(�4E��)��.�����I�.��ce.H�\h���۷����$[���+ٔ,�DŻ'�4�)����x|ԛ
0�y�x�K=�Snd�r��GZ>&\c<{�=cI!�6`���{W<A�x0�݌��� ���B�a
z���<�6������%
c�*\89�����p|�Aú��j�}��W��WJ��Q�O�K6�P���-�9<e�ړKe������EC<�핧<c&����,�-D���wơ���i�7��7w�M����K^%C�Q�*L��Z�o#�qCy��������H��j#M�W�J���X�<��ۯS��Ws��b����݌I%a���?yVC�z��؂�P�ua;�V�P�$_
�y�p�?9��dI~\ҹ�j���ۙ+T�P��PER��X�sl߼<��M�
��Z�;�K�N��
)I�	D*�7`.�����22"!q��bw�܆D��
r�7�f�qY¤HU�����lSn� 3Σ-�Q�d��%�M�rG`ƻ�NA4F0�8�%����r�����ֹ�Z���bŇ���1=x�F>��P��c�`͑6%�V�j��vf��Eg�{�LO���AZvW�c��p�o/�:P���0�1A{?H��#+q�6@NyL�0U�X0|��zUPõ����=�
�B�65�b`�R�#��y�ʢ.\]g�>�B���"�p��n���@�vu~X
���kQ٭Yɑ�&��Rh�����8#���B8F�&���Lwޒ�E���=��LJ��G;�=H�8B*����>w��O֚���4I��k��.SA�������7�n�Û���)���`�~�����reryεh|�>�(��U*�̭�g3 �ɲ3]��\Al��^�&ᘟ�/�]+a�Z�GLb�Gv!�8N���Z֨�o�P�c��YG'���Cf.�$�@����~2��u����H+U6XD1X�����@�HP���(n���0��
m7�N�t���O��I���I�9<�&���3�rSoԠc"w�`�1+rv�C���K�HwvEy���G���8��Y�,��7!��������y��??��'�@3��%��;O�9��4�D}}2^g�j���U�gk�!Ϩ�3��n�R�MC�y��Kތ'�R��vZ��y��x���q-�ک�@�|B����$>�@���ў[о[~L�o���[��������QO�f��eU�r��1>��Zw��#cӢ�!��yҠ����i���H��5˛����ld�3EQ%�>�{��=\����(�U�f��*v��B�G��_\�3�|Id.m���������+��w�ӊ��ǝ��R��������\)�ɒ �ŵIL�XM�У�<���a��/��=&�sf���Qg�
�ρ@u/���\����QM%T���͗b�b`�-������ir�]�!XP��_[a	DQ�ǋ���t�E ������攒�&A���(IDջ,��I�P`����o�M�ȬM����l�Y�V���*��:������(�y#eU��+v&�ꠄ�G(�$�/t^���xE�n�(�℟�� 	�����H��|fYH��O��S���9�&�E�F~�l?w�u�<n��T�����!ɼoF-�S8L)k)���wf���p���
��L�4V�#P�`�w��1�m�rK��3�G@�&7N��Ƌ,>��瓷J�aF�%ѣ��4��uP��+y�p&�8�(eO� H5/��@�'����b�o��{�)�b�*�y7
�z!KO[��?4Z,z?�/a���+MD�.kt�v93�Wn�)^���!mtCd�T2� 	._[��-��˔�����)ك-+�8�ȉ��v�9��Q����x9>o m�����as�w�dK�v9�::��*}��r�$�N:X��j�S�,�Z�e��GNqd�|ټ̈́������Y-b9�:C��,�%tO�A��n[��N{K��<6g� z}�B��6�R�w*��ǲ&�Y����t��b%�;ߡ=Ea/0��צ"���=���m��ِk�dP����Æ|9�	`�kGR���Ng`�Of5��M��F}��g���x��=���.���aD����P�]d��}����{[�%�f;)2���K�b�Ul9���b�fbD�?��t��=15U�zA��-A���1DXR��7::�Hˣ��yy��"��f��ZZUM��gH��el�E�Kl�g�ҀY�ż���ڙ5�J#�+�Y�nu�,�wfP$�Lz>=��*)�ЯF ��:	�=F�w�`��I��}�l���7A�qF�wR8zd=x#��Ŋ��E� ���������}ખM�����Y���b%����e�f�6q�L���Ѿ:Z�ىa~���VU��w.eE�>��y�4&�9y�cO��0ᶝ�;��D%�3!%K"����(�����E�т�������8R����;�Z�џkJ"��)*���}Uv�i����K�W0�|~Ds�B�rySēnV�Xk�3�C����לN��{q���j�~�P��}$O������#*-}�+������Sh�}�a]9&j �*U�ֆ*�v7@\7T����?�W������|u#O�������uE4�� x��Ol�3t�
�/�Ц�~��o��$��P���=�*,��Q��-V���WqKx����#��3��c��X7����#E������=�"�G�/�C�Xr>��#n��դ���6�t;n��1��=9�F�8�eV�|z�b��l0����"
|���C5�Y�zŇ���_������ �y���@j&>�iMR���X����ƚJ��a�7i!�JtT��>g�4^ּlc������>���EK*ߧr&�	���V��g�Pe��U��|�a���37#�<\q�I^N�E��Q_c=O�áv�Z�'�5��4��j���!���7Xů��9��|͟�V��A�4�Hv�7g��X����~SS�t,Z�E|M�T�ަ@�lA"-���<��jϵJ�z�'���þ$��~Tƽ(�>;�IKNlqYQ�6���p�=���Jd�	�R[o��Zz[F#�tK�U�u�(^��n���eb�9�>��m��V��뢗���4��fP�Z���QM�"Ѽl;mm����~@�ߣ��O �p��XR*]��|�&n>��/>$pZ�$$�	�f-��9������׎�����%5����D��$��_����pp���j;$W�PۢkvNt6DmD��{�K�E�����Z��#���@r��LK�b����"v��rL*��Z���(��������7��!v�a��u��9֬y8�7y��\�=4�B����z[�!�_� ��>��������!^�0qyt ���2�$'bY�������	�]�����gq�����M���� ���A.3���S���ӏV=��G�#)�`բ��͞��d���W���T@p����,�.lT�.F�>}�3�Ju���l��f!"(�4���v�E�g,
�azo��7�k���p��=�z.5�a�Mʩ��[��Ѡ��GA�u�;~�09�1��=���Đ�Qk��#lrS)p��e��H:��)��(�$���(@�"w���kkUd��Uh M�I�f5�Q&�dGA���Bh���p��㑮�W�Wdːu�eU���������$V�]c�'�HRP��b��'<:ϋ�� �4��W��& ������<6���̤���0�N[��="���E�ψG�A��r�l��5%~V���ҫD��M:���^c���P��]
��N��]4�gt��W?g�R:Į{�lw��UQ�E-��U�L� �(��YS�(�u����
���,�$�:�K�YZ���-(��+����믽ZGjB��M9WaG�#�>�a���>Я�Qǐ��D���dk���^�#-?�O��I֌�[|�#R
��P�t�[��d�F�����3n�`�0�Y,�¶"��
�m�����+X	"�Y>:�na(1��?(z�5/��~1��#g���αaC@k�(��d̈u�R%g)Up��S��{����b�Y?,�Vψ�I�}vKHїc�~Vk��i긙����*抣��e�������j:�B��Z4
Լ��5�6?�?AY-�KI��J0{����~���t�m�V��"㗮��;��r�v5�$�<F����d��6�����3���@wI���V�V0{�K-��i�-��:�x�τSG�]��RR�9�d�sEO�����Q�ߺ�p��ч��(-׃�x;ª�	��a�O��5(��)�*ƣco@w���=�:��=~�o��Px�(�LW�A\�>�Γ���l���*w�..4���^T�nMb~H�DDi�9!���c���G���odHugI���c��(쮐���'�i�4�q�:���J�=�iS�z�Uޞg?��ﯓ�d�,ul%Cr��N	������Cs�g���x�ͧeӰ٦"�m�*�ZҌ,��̚���J��},_{-�2�oBμ$�m:��e��}�ԃ�<��/Rl�P��^�n�{�v%���$�d�S#���u��ZA��
f�s�+����wsg�ۥ�����7��X�\r�1<>l���2��Fr7ɘ4��1��G浿�0��Q��`ʟ��=$��
����^���E�ʈ~�c�Ӂ���^4�Gp���q�^yPR.��GfR������}�����6B9���:�����%��R�r�e�ţ�-�G僮��~TmP�+�V�	k�NloV	�R��}���ƿ�n�QEf	Rak=��K�F���Z���t6��x�Ń��,��>R���j�T��C4�p�= l/���>;��-G5��F��,/��%�/�M�W
��V��q�D�݌�n q4끝���SA����:��)I��M5�k����m�(ص����RA�g�Lb����m�4�!�ieR��	msw=�S7���It���?�u��RkcW�"�֠�<��c�#��*8�xׄUaW�-�2�}��F�b�Y嘷Ƣ5�8�hr��Ԗ�_���C�.�⤽�~�`b�����7Uy��^�|	�T��G�0��V�:A<!���d �tǬ�����a�\����n��M�e~Õ\YA���y���#i�~�6��B�hy�ƺ�f��������G�~Uk�柕������'Y�Y���ۮԻ���K*��v]�k�m
�׍~�K���.u&��[��_H]&<�2F͠���݁]���.��*�ۣ����l9XO��bP�L��S�:���b�g]���B�����N�"�p�}&6p$m��D�3(/߶��/���\�_YV̰��k�f�����R®���&���:��AA�s�]D�L�7�7oGޡ��z�bw�͒f\�l�r:��[G���n��	K�-�W��1�����p��������?.Q�x���򯍤U��cil�+�2�@�-����	N9Cn�8Oum;A"D����F6�s`'J?��Z�I9��%��f��ۺwȅ�vpH���a㹔0�`�	a ��oV�v?��R�=�UeU��>��~�X���j���3zj��0�3��*g�H�)�2��D�s���ӓ��6#��V<���\�ڴ�N�љ���m�fW0PMy`�k]D���V��+�7�1s`�k���C W�HUDW�K���+��`�"�w�,��f��}h��vD�;h�*�P�Q���"M2wS�=,�l�;���۳�\����~M�ӕ=�D��'5��L׏���˂��l��	��-b%�sɓb/�n��NO�bFJ�1%��$	���U	��G#B)�T	�m�C2s��veʗ��Q��0�H	G�H��� U����5�|_A��u�/�Y�4#�F+p������R��æ�w�ģ|]ױXuh���b�^ntav��I�.x9�	�/�t@�������x
��9�a�yU)g�,VR05�b܁#6����ɳAX�'���+��,�S�	M�L�<���vJ��z!L��ۡ�1�r�f"�a�	�1.�hya'L%�<b1_ERPy�_�p�ؘ�g�"6k��t[����$>?�$����ԑ��Ix��0hY�c�o�'��5J��bf\kz�&}h�¤�#��1P˯Rg7'��� ��A�|���8���P�w����'7X���w+s�E�p��S$붒J�xX��pٳ�oO�B�h{�3L6*Y�S�b%��So��>�~_����I��m�;D�3&@L.>�&�\����d`�op^��@'�sM��d��C ��{[�0���L�D�q����&q�*���'S�@��G���_ �{�P.�[T��H��9OM��?����u�������;O�m��J�S�S��gd��j"��!������Y���:�S|�&v-���=�<l�������.����J��������kJ���^ӱ3����76-�Zg�F�Q��!� �S"���Zz����z�n��Y���5���q��V���f����w����OU���&mr)������Ȝ=���~�x�)Õ7�*�q'�C�C��!ov�(�n�E�9Ӽ,�ut�%�z�}�}�уi�:9��_�������N��?�T�~�cH�<H����v��1n��J.�{����RI�Oi{��91����&}����º-X!QK�=騵�B|���Z�쳸�H[a�a
ں˱�/��k\(���Ĩ8ā*��텺|c�`ȘY�(��MH����̮��"�m�����EY�\��(�W��)ḳ��2v��C^Y�P��ٳ��"�KW	�M���� �4��F���E�s����am{o��J�����}�+�h6z��]����D�W�����ǐ�g�vaF�=����4;�'��V.		y�P#$)=;\#??�EA�̚��^Re���E���t�4�0]�K�_x�*�c�]�D�n�v$��R�6tT]���VQ������.��1�>����aZ���c�Ә��y����g�c��D���	�w��9��PP������T+L�=�	��ºu^j�;�'��:�mȞXf�w܆lp���a��,M+4�S-����6�L���$��͖��U��	�S?�.$&x$�LIo�����^���4ޡ��l�7vh�ÈXd[�긐�
k��ӑe�,t!�[%r$/E
{���E5�	�&&�Xv9���&�xKE����!�k�����f��Br�+���-��&�]օٍ=Ko	�L���H����Fiwo���}��<kx�!���Q{�}-��yCLlT�"��������_���s*�BЭS���u�k���i���
�j\���IGv�h�5Rf��k�������2� �n:sQ���_b:���/^YL��.���p!5r|/�g��8�g9��B�t������`��Gǝ���Tj�G�N�����
��\�F��M�@'p��G(����]�W ��Vo��y�A��KS���y���l�c�t�
+l���^G����Â�p��=�\0#�����R�P2��{�$�oq@}8.�1�s��/w�#�-Tt}El�5,ʩA������>��l�����tK$Z�h����i��I�rv�QT5��`�,��1�g�����*�����Y(Uۚc�o���Q��9�l�vyl8�~0G�Z�UE��jz8�Bj�������4�h�DUcX%a��	�x�5��} O1�P�#��3��8�|���N��ÄZ�ԛ]-���y�\^����ss"�A��$^C7dT1�ȭ��Z/{0�ӌ�5(���5��Q�5�A������ϥ��1��YY�☫�M~T·&�k�SI{��5����E��;��:#��r��'�8�}fa=���32v ��w�yu���E�Q��n�0�؝i���`x�%��g��R�+[�t�e��p��X��7��`W$@{>W�z���uFT�%�Z��F#��ۆ;���/w�tS#1hfN�%�Q����r&� ��F�'�̐�Z�)�FH�k֐s�������]/�=���/�����j�H��7U�	��[�s}��W|�V����?��h8r�0��>��<�I�GTl�x-�lx3��I�� 7#��{����zh�M[ᬂB��}=��=<e7D>}k�#�l<TOk�n:#��>���]:����j�p\ߥ8���R�{���]����$k���B[�D֤�:��	x0�QFvų����`�����/�̍�9�RfG�S
���b�7�ϭu=�/BL���~�z�#������֌�?��)iK������
?�
j b!�g��
V�E�5�(��	���@@���@U��$x��fi�;�I�'� ��K%�����l���3���E�ͭ���K��O�;�:)a`�"T��c!�B�(P�;J�3��5��<�ۺRֺ�g[���Ay� Fu�ρh�	���ܒ�O���Rf;E�G�z���\2��"�,_u}�fj�6"Z�<L��|.
��<�5a>����_��x`�-g�AQ<�bq����|��c���Y���3�e�E�r5o��Mߊ�zef���wA޷s�5�����0�-��䐵N���0W����+��?j�"��l�;���%9�Yr e��@�󖜠�����[�����8^J���\�$\���:�f�JF�������m�>a�Ն�=rn��b����	�^���K�H�j��$���'T������7AcL3S}k��bM���x�azl�yk�k :[`�ʷ��LpG�*�Gp����[�:�S������@W��m�"�٬r�2NE��P� ��p(DM|�T�XVZA�$�[�LnC�C�Xt,^yt�Ū�`W
q���d+�q�9؄x��p96�O֘p�v��C�;Z����$=��Vk�wE�>��a�b�5T�f2:�.sMa|/���<N�E[�K��p�<����P�KH��'	�D�����&RKS�/)��uc�|�gmNcU��? "g͡�R�RC�ئt���-��
N���eَʋQ�4��}D�RTVHX^��R��{銞]�,wY:��ֲ�{���1�Ք�{�����#u0ǆg�W��\?`qo?v;�ϴ3(�����L�ʅ���w4���-�� �8=D��t]A�)��e���_���^ZI*�Elt �����K�8EF��X�K��3p(K�RZX��48Q���]��bTd�"��M,}�Ph+��&��?��#���6�
���jkZ*�z��R�Rە�]p�J�?E=��Z�f�Ma���p�[��g���?��q<�m����w=8�eL��N������K�5�cj�1v��Noi5QJ9��_u!̛X���g�S�H

�NX8�=]�s7O�M
�f�t$S}D_�X�{'� �5�\DB(���D̥��ۿ����R��Y�fnb����DYt4۽qkC�C[��Ǽe��ʌ�u� ���z!�$��'!�P�0���.�,ʰf�9�܀(����ڜ �mc�)+���Ը.\�>��ί�s*Ԙm�8`4��s]�; /����s�k��)[] �2L�XN#�N�b5Z��x�e�[��u=���N��Õ६��i#����&�v8�������\�y@�k��G6����䉱j��8J�\��侒#V�e��mR�@1�*5U�V2�Z����������)��~i�(�>�?B�.݋!]��kG�j�o�!�`Q������]�eT-�n�������J��Z�����U��4�x�<���sV`l]��UNzZ���g��{�(K.�Uvz���_L�\��)Bb �w�!��ա����s��b���CI%b&���O��tP~���ʹ��U�@���	}]#@	1�&m/jN���_�_���Wy�=��T#�q1�c>NI&8���@)�մ�
�E��H��fD�jI�#ݨl]L�[�Cˆj;��g�[��,RX89d��kA7U�������C@�Q~g7&ЌCO5�}%���^
�u��$g��&���u�N�|�w�r����5���~��M�	������X�0)a�4(�D���{���l����Q�A/�
���~%��P����٬>����NY"a��f�4�Е�T��� �c��~$��J���l&�o#�Y�F��_$eщǈ/�J;g6}OuV_'@��no��{j�fg�i��^Zp*2n7z�e|��d��Js�� �������T,�|N��1jՎ�R8'R)��X��߽�l�.��G�E�-���������2Ի�sMq&ȧ��� ��;cZ�6Ú�lS%�d8C��,1�I�T��t�_���fH8�c9~֎q�z�ǜ2#|ARA��n�Ko�Z�q�=��������70u;�H����ȯ�*�A���B�2���7򀰢�m�p��S��3�+���b�UN�Ve�]<�>h�g�뱫Y�DD�20�}e{=�a�	p�IWڒ�{��g����+�����;ț|� �-4L|�RN|��^MmX~K��F��*|9I%
<�g��$��Eb��.fR;?lY��O����e�~��p�'.8�z�W8H��7���R=G���10n�f��э�� �_3ēa�Xo%P\�.&`O�����yh�����B`�S7�9X��/	��t��uv�?�(�dÁ\��_6�W��w�j7,IG��iFe�h�x��G��*i�a�ݔ^=�h�fj6Zf�YE�C��zP0�����fH5�?B�A��@/�ԥe1EwQsn�]l�����BV�������~��͂��zwa�~��_�T�[��40R��������q���z�����*���>N���-�������^��kui��(kZR����qx�7���&$	,�vK�!��#b�x�<�1������4�������\_�6�����Ze?�*�6˫�c'u�Y��D
�r�sF-�N�)���*U�2�jr�ax`��({M�q^��[�pY�GC�`�����z�/�ݽoc�䕍+�ߝ�N#<�	�0�e����I�(���	p�C�?1��^|� ��"�B�]Z��x�c��YIÏܧ��I�ա�0�"���p��>�4�K�fF�m#�Sp�d�Z�:��<"�E�u� L��eD���<�L[ �_^\����Y͛wZ���hr�m4�f٤�d��J�4��������� v�0�[5����2��L(y����t.�/>t�3�ɯY,�x�o��GW�7{z>п� �y��Pu���Fi�+�U)U=�<Rd+�T��_!���X�X�FEl�«8�M��fu��ܢ�0Q�t�Y��b9ݢ]{IJ
�t�W�F�6� �U�=R-�p_��x�tӦ^:��4��2
5�O>VhB��6KVe\�s���.��5�?�{�pK�ѝ�;G�Ȕ?����+Ѱ�5���!ΉOFP鉎����� I���0�>��qJDtQ]ͺ��&�fO�AW�F v7sę��9�1k{F�dWjs"�| �p;��w.�`aUI-�2��R�$ZĠ)�7K�6�����y#�$�?����5�H��G,U�=Zc��D��!�������O7�j#�`�w6�SIQno2|c���8��e����0����\����:{�p���^ቔ|��?���B�c�ӑ���7Uo����HJM��S�}p���<�E��hfR�5E���v��d���o��U��>�jP���n���>���8f^�x��.TF8 �H�N_ �"t"�E4��+g �����׿�
�)g�S{U)oƸ�Z��Zr�>���W:��~/��ކۚJ˼H&����6$?��^�%�iȬ�H��_Da�5Z]�k��tժL���Q�I�&�h��fG��+S���c�z�,��B:ҋ�N�B�)zI������zj<-��y��;]��������"�[��̞]v��4�Y9��Ծ�ȭ�}���ru���<��A'%'h�g`b⳼�P��;��������|@(I�/#7�Z��%��T�?���U��I��/xPM�;�Ȍ
-N�7�
Zh�3��
}~�Ze����J�-|T��WI9-gvvy�@��
O���(y�E��Y*���(jC��G���m��u9B�����t�i��C�ee�����\�!��ɖc��Wv�ή2����ޭ��27��nC�#��Y?��9��[�	-$���$nm˵w[���S�?g�bb�@O�����$�^�x�:�O��������9E���R��D�T�Olx�|K���h?7v�2"��;O����&����o�S^�w+��;�aW˰Q�D������b�(_�2��:̿D���G!!�|����/}��\,�e�B)�����a��u�1�k��f�2cMؗ�'�<\P ����t*D�P�+��8�i����Q�
@4E���pE.޲�x��;ָ��y n�T�0Z��a�"P/�M���i
$A�����2�M�9��ǎ��ry��ϳ�D�� "8��e�+=1�f�d${�'��#��� �?��w�)āa�}|yF��Գs�:�lD�T�cg��/#��"�(���z��u���.�.=m\��C�h��U��z�(Gl���^̋��i�$��E��2�l��a}b%
�W^f�����1�d�M\8����&8�������X��W~���r3&C�M^9�m�n�F�H���	n�UO��Fe��$5��Xo�}H�Hנ:���.��j@j���JJ'�VR����%�'N�[�*A�W-�}L����l7����?oS-�s�✗�*� �-�+V=�)V"�|�D=�J}�	l{}ň*͌RaN'��^d�����g�_�*�B��V��L,Z�<r���_<�\�A�A� �D��do#g��q�� cѺ�4^�Xwz���1�������<���G�7R����W3&��uS#��~~�o��ӈ@2��~��'u��ϯ?�9[�O[M�'ơ��+���
V���H� k�bZ����[P=2 �T��TOU�S��]�^w�&��+}����
O����i+���m�yT��ӵ��8�� ���4K��5l�*dZIm�k�M���`*rYΈ��3M�?����p��Z���h2M��.K�zV��d/g�$K��r4\=f���h�kQ'RD���N�_fLv����q�?ط 誧?+Xw�{e��+�F������\���	N앞��5���3R������E�� �,-I^]^G��&t2���^�q#�A٬I��?��Or=|�L��
����eJC� Hr�(��;hߒ<�7���¤
�>c
����mפnb٦'���=��f#�f§{<��h$�����c��_��O�}xT�k6ޢN"굣�A*Z9$[�p��tx �9mp�۟�$�?s�����E�.ͤl�z}K�C�x��,e�2n
Ή�D����y$�}W"��MYF=�7����\f�	���⧷�7�d��F@z��J��i�T�nFJ�9 qO�Qy!}}iK�M�=�ӄ���c�r%�1~(@p�P�_h�3��kâ�C��chE�L�0�fy�7����Fu^3�kWX����AXƥ8�|q��4?������[�c����S�ɭ�&% |~�a<��R\.�9�+��&��2Wn�.�@��,*� #����)�u���$նE�=�>|�p>v�p���G�|;�#���T"ói�[�m/�	���h�ɿ�>�Nq�Eh^a��y���;��L3|�_8>��.
t�j�s�xf7���G{o(x�Чv�3e�ƞ�˘_i��H�L�:��C���J5_@}�ډRB�|�_�&���GZΏ�+b "�NX�-�V�X�D��k��*���fb���ȘIs��'P���-�֕������VA���3!/	�dmh�P���ZG�h$�A
�&z�ұ�!�78\�h?V�P7�q��f|�H�Y�f���q�A)Mlز���b]|����V|A۶�t��?�6����Om�����Pt�Z�+;��Kr{E�c�I�iwR��j�|>���Q��p�=�w�r��l0"Ii��U(��GE7+�o�������Œ�!$�j>�\��x'r >`�I5�S/z���n�K4�����23t�p1�s��C��WT�nW���$l=��wG��UZl�h��xw���Q��Ɔ*x��AK,|���#�Dyw�o�Σ����>uK��aV��榎I��ĵ��_��T)���������u��!_A����Uq���I��#Ɓd|O����Y���y���6����ٮo|�`�)�jQ���+4�?�d�|��(���у���ևK�?�Q��*F��&n����U����B�k�@!��U?J���]�ϭ�v\s)o�
V,���I���"!"��du&�eO/x0����%*tP�:����~�+�J��#�ң��� �������i_>���a]�� ]�QЈ��x9W�3 �����!7͗X?�����h�̑q -���"�Q�{���藒S.{VF�`P����*͑�S�#�b+y��P*���@�4<��!�c�Q�����>?:B��:زK:Gl ,���iG���Yh�"wW��O�SC)��6G|���y�_�>3��@����<?ĭMqb��5�gn�IXCw������j�a)�G�ϟ ��8���-�+�]LCOK�?��N��Gc�,)Ы.-sߖ�;�E�ߡ���g�86��b����$b�?�orxȎ�§�o�kd�9�N�`�q�3NW�m�u^����+�	'֮�n����%�Y�TSF~��%J��|nc��O�j����ov��1H-W/*7e=�,l�Uޮ��́�ӟ��>J�^�|�V˨$"�2Y��i�w�Gqo�`J�z]���Z�Ț���rŌL���T���$��"@�r��Z��q`�s�c�;�r�+>�m���|z��6a��-���?e.XG�6���:"�YC&�$R ľb��u�)�G��T�;YY�$��{^m����8����1}��=�S���Lx��w]���g� J��!�x��5{>��e(����Y�`�saM��L藄���k�c��%ݔT�l�+�Y�Kʒ(�E G�����_h:lA��%O����C���/a*�7�\�2��gv-	���&��.j��	�Påo�x���Lj}�+��Dn�M�Y������v̳�2��d?�w�=tΌ� G֔��*s�H�;���X��n����HMq��6�TA�(
I9<�0��$��=*��{��vP�L�:��0:�+`���rG[-W/�r�]�P�"�����ϔH	��u�h�e�
�:�Ǹ��"͢���f�<C.>�v��cW5t�[e�fmT����$�r�\�&T»`����Ћ��k��5�y[).���z!���rJ�޽:���‐n}��3�\����^���z�|�{����!�D�9иi��9��l��� �|{�����^����;���ٵ.�Jw�r�+w�d�΁�/c䨣Ǔ�,��H�4�f���͒���'{�t�����ɯ̾n�z6�|��k���&�#��i��Xo�|������W�-c��م0�)ʭ�S����!�gp,�)�|
��:����m��bnE�@Ҹ���δֿ��ڞQb�Ђǰ��w�=
�)^��0�]F�<AiFت�}]�I�� ;̭)$�F�χ����phJC�e'�ᕳ�րH��լeû�_IQr��Ÿs7�S�
!����B���2��վ��@M�D+:d�#U�{y���ˊ�.b�Pt�Z�F2я�w��7��xb6و:����d{��ŧ*�j]C� 1��E�D|4� �G=��08�;ϙ�=#S F�����1Z�o5!"�
���:�<F|��0!����)�s�8��T;;܅���b��W�B|кoBq[,��t�=�/���%g�e �V�l�FA�T�0��R6�}�hy��,�b�yO]e�:.%�aw��X�"<�K�	�LyN����t�W'N����ݔS�d���/2G�+���e��z5B�%S�}E�Ψb�����F����xt�ˠ��l�� �kK���FS���)�Ҭ~�<U]�+�uˁ��V`�~��U��g�(R����G1�����l��h&�>6��k@�HF3�P���U$R�~�x�N�vc�Pa���t�j�X��C��ƣ�������	Қ꣦����.� �WVP㍣6��=/�VP�Z��C[rRvٯ��\��� E$e�>��x)��~��z�)�W����"��$�(7vݏ��)o�߹�7���c@�\����?{E������)��A^��z%
 �2��i���L�`�Ƿ�b?&,�OcBf�^��kU%�8��V�_mO�����Ai%�.]P�8��.�"�/ Z82��_��w/Ծ��K��X��o���a2��\���:EJ���.��6͌�q1�W�ťt�ܵ|�~ x�L"�V�{�d۽��?�$o��9�Hpk���dG>mY� C�����C$��i��8����H��2`.�Š��yR����;+�~T�5-G_��]�;^��{�c����F27՚��6u���/��j��Z(�!�U��4e��E�~�MN��b�����M/V����& �;Iz�~c	�`+0 ��w�1uP|t\�sc���+#����o_3"�C☪�qaz�i��I�t�|H~=��'}�^����~{8�\��&�}����~�,�<����d�����`t~�h�nQ� r3����¹�u6���a���7�[<T\��������������v%[/[u��afj8j��E��
���shmBD��dC��f���Դ�떆8ӽ�ׯ{�#m%b��i��(g�|Mn����.RmT`���3z����Q�}eÅy�0���!�c#�f�l<���ii0T�"0�x66��>�d�>�Q�A�"���eդ5�K��]xM`��R��zbz�I!����F����?��̈́>�*c�͡H��,���>n
��$�Ș�k֔>�l�20����e��"�9���E�h���J��:��V91�g�8{�|�Р�?8�����37:��+�1�4�VF[`2�L|������A��>1):Vq$,N��s���Xl䫯���H�Q�W����
A�������;b�
�6�O\�+-�wq5%�~G6h��������Jm(6)7�r����ju%��Թ) Ԟ0V��ϥ��Œ~�+[\B��gGD�����l���=l�K[p~:�b�k7W:\"�>�}�T�������x6�a��5�t��譚~N����W����i<�abCt�"sǊ�P��/�kM�$�	U�1��}8���5A��^����U�g�ϋٮLb�0Z�^�&��X˒pyF����ޒoc�����1��ǢQ�ue�F�.�_&5�-��������j���>N�ve��w�(%���L�(��Z���)�AlAXЖÂA��:T)G�T�S���w�����臬Zm�	������#l!��� 	
��R��&WKW:X�5:+�t�%�Q�k��1B9*����b~���[��N��n#�c�����E2��y�jJ�G�b��Mh=t���h۴�D�_��ˉ��&�z���֑
�{!7RE�[>�I��!BE�˩KN&������UTyM��H����roT2l$}@�)�W%Դ~Y�{���\/��Ț?D��[x�Y�q|j�!a{�̓���6��a&{�{ǜ�"c=�������ٻy(�kB(�-��o�0f�mt@�uǦwL�[����d"�"�a\[T�k�h����J*`p�ݼ[0,Q'�W�j\�ڍ�
��4E�a��.P��'/v��y���RT͘Q�Q"_�#c���S�Z僥�GW��%�B�|wU�#��I�;z��2�Mb���z����~������v��=^�
��P�}8� �-;��p�c����XS8{����	���U��ѣ�L�"$n̞�\��-lg�M6��~�	X�.7�@��Yн^K]nk1J����MÂxDo+]k�ӠJ�����0��=-�7�ɩqԎ��Q���ݤ#Ԕb���L���++���%�O��,v�SKr�W�d@Z�0H-_X?se���_���10x�� ��� �#_���q�~e*��Wh3$u��bјے����h2����b��(�g;��Y��H��i��]ŭo���2fO�5W"]`hH嬃�@K�[ �d!Cs/$4 �Nw>v����=q��I.���ޱw��#/n�O9s� Q��^WTC������\������IZAC�*�{��A �Č[�5H66֭v��<5��a��o�b	��� ڇ�2!����wp��%7���ɲ}��[�]��A �C���m�*w�'��Y˻���a�An]���/��hЅ!�|&�u�!\��o�*�eC��I���dG+;S����)}�r�<��|�R���9�����kn{j�̷t�i��>���/l�'I�Ԍ@A#ш2���4Dt�؉y�N(�������~�4z�/m����&��P
ě?ϱv���:�v��b=0��	f��'���er��.p�8�0�J@�����H/*d�"H���?���m�1�7�v��^L�Si��M�g����%lt˕N��+��-\T���c/�.�y�y_6U��)�.@/L����xt�����G�x�e*@�w�<���Ƌ�8�J/��O��Ԋ�������d�qn�"��eY^���x�N��E3V5���j��?�(.�1ca�6�4s�8KI���W8Ix��ͽ��xo>HV�H�G�v�࿍>־�}���71� $+��&�k���P$!�ʜ���`_c	w�֬3=���Cd{���ʊ�LP`CC6ruEn��J"����Wt�[y�.��I�wi���~I�-k�?��z�g�nR��8��<�2y�����v�L�e��<Ւ��T���B$I�}���6,T[���ϳ�b4�An.���?g�
ɇ>[��	͆�>R&ﻵ��������de{�(�>�>��9�I$.�5��5e�
���F�mp�s����$	�y�F�v֖(����kK�C�<#jX"���w���{��/!�\����'L�to':Z`��m���6��"��8�>��}�y�z�W�?�����b�P�������h] ��hO/`(����7g�>܂uW�h�϶�h�^����G���2���Q�s�	�8�Ho�k��P��hݚ���A�-
$�˲ǋ����<�y'()6]�xWK�R~7�arZ_���9��T�h���[[(B3ǌqW�����t��1T�ki ���������Ka+j�9T(�B"]���� �H�h,��P����i-B9g�䇁n��>!�^����O�N)���n4G��^�@F��[��=��-B���	�<�6"�`�U�}�����i2sb՚�|�>o��F�	0e#�s\]SF	.��zB7a�����:�J��rO�2��p!`�p)\��d�G��Ƀ!KH��?Ә����ޏ��80a^-���M�=-Y�`�o$0�`�hHm�%W��;��0�7`9���<��{p#��y�U����=�ŌI��V&��QGr۸�T-��wnZ  .ө�J\r�A`݁B���n��<��P56�x�� E�u"��w3�v�ߚ;�A%�ɗ=���\� R	&�|MJS��~p�ˑ\�ݦ�1!�������!�+������z>��W�B�M\.q!Y-.gX�����������'>�q�N���p'�'�s�*� ��1o�h��Yt08ɵy��U&ǲ�_3#Ҧ�$֫&��%�'JN�W%_�Ĳ-G>4���s�?�������M�`B�0���AL%���(�k��6E�8���xӓ���}ҁ�hW;û��W"�*����߲�G��s[�a�~�U�3��}+�q4�������(�A��ٵOF�]]'����yT�s��s520�g�|�.��\���B�����^�-��U�#A)�82�Iǒ�Y�F�w�piH#��%�T����������Qb]� ݹI��M���������C���j�nި��ȝ�0�3Ye�ԝY���v�~�@�PDđ��5�!,�6�2��)��X+�W���W`I���n�G�	�{1�Vh�N���/X]�BZ��x"��@�]��1�3�r>��AI+f���e)���$�yD6ZAM��%�oR�r���X��7.~��E�����u�yN�XYf�|p���"�#YӢqzq�"�c_�Z1��#ˋ���B��*n���r���F��:�qY��R��� ���2�woT�*�P��y>n����U���Ԃ0흄��<{�����{}g8H��fަ����f���t��?zW�RҤ�t�z�x��o�`m���ss�D��W�,�Mh���=���$8ߎ�-��{������>d�� �_�~H
�Je���� 6�V/;�Y�T��|[^��@rS>�<�F���4�v\�1�$�1�H�;�Q�#�CHݶ1��7���`��w=�)|��#@����@�� �BL�Jo#�����#�Iŋ"�,J�p���u9��O�T� �	�����$Ϩ�Ѓ$�����
��aݾ�[Ӈ��O��^|qC���J��o�dQ0t	�������@6�D�H���,(Ӟ;^��*2 �XQ�~�U&�����U�R���a���S���Y�_E�Pi�y�P婘g�'S���*G%��QZ�"*��}&�X�Z�����ʋ>���ؘ|�ʹ��[F�6�P���=�"�܅E�7U��&�&a�6�g=��~V�I]���!�k@���IC��l k�(�^U��W���~�X�
���nQH�������.Ί�(����3*L���辒vD������;
aQ4��a0;W8�Y����L��W�e�W ث�DN��
�j�V�5��1��Vv��m��\�������<�2������_�7c1��1��Hx	':P������Z0���K�c�3ʉ�u�b<���8���y���Y�ˁF�^gs<`��:�cv�P}�M�
&$�	�,P{w~l������!��})֟6j����
��6�|�t�9NTY�T����ZU�#'8��n�����ސ��P@u��?/:��ځ��`��@֨u�1/�檓��[��G�������R�L:�0�E�y����^lO����@�2)�(ݥa����x2Pkp
!�5����\F�J��'b���Ǝ�C��O�&�균��;�;h~��%f��2�V[n���JO��[��J��F�K�+S�r% M)8`�͌{�b<��Q3%���zXG�XŜ�C��aS
�P������%��k�Ad�+�T��GX|��B�����)�f�ݮ:Wf*�`�FP�P˹e�[%�$g�Az��E�5�Y� ���G��O����i:e���.�$��b�C��h�`e
�H�>[�F�wg�׶ }������^:F!#� ���'_����4/4���Ӟ�v,�L��,�a���o�X��ґB�`N��/��DfI�e~U�	�OG`[��qZ����T���@��*�PY�[��D�S�8��Rd&l1>�vB�K��޴"��-�R�Va'�A��+ꩥQW�)�	ot��Us+i�Z�Y{`:��£�F��--����1+~��E�����'��s�;Ğ�9�PŁ��Y�yk�u�s�q>vc��H%�!���;��
�K&��m�h	c2��Gue�*d�L�f��<��0�̢&]d2��n-J"�/30�v��۞yX�"�B5���x�GJ��-�[N�ܘ4�%��lE��Jh їG2[ψ��>W�yC����9�Dzn�p�)^���N?�V al΁�v $�.haR��CAVøҩ(�"'��y�7�t��NI�
�r(���2\"�,�UVv��������5�ky�S�!8�v�-��I�l�N��l����#�Q~���t��g�5ԐgM��̧%���`�f�@���I�6��m�q��ECJǫp��}|��4����_��A���S_[}�ɤ��1���4~�k�0b�j�N�}��ԿAH�m .?��s��%��=�wʅ����eh�i���jy4h0�h���_E�̄�.�@-��}KPU�
&֡5���ZƑ��`o�����X��q�?'�T�*���8� �I��V��څ'E��{I�8�:���osg�Q�߲
]	{�p�~JY8����AD^]9��6e,���q�/�TH.��(-DP��ŕ�	bd�-�˺t5��s�-�3%��]lJ�,�zE��@cm�~�8�e"���$zt4�Ye�����h���A�z�ǳ��P2�%w�/&3m���F����O��y���?��.raX��,T�P�b�������A�G4.�C�K��`� @�ז�n���s�]�I]��^���G��&�nf�"K�N>�'���r�Š�����q��,�BoUɲ���y'�p9q�2�����g��`�2N��Y��5�F�YpŃ���<dNȅQ�[X��/a��c�m$���	��N�w��w�$��27��A��ù��Guȉ����\�7��qSWGǡu�����6aB��$�@aB/6/W���У^}+I�ᎼY������k��m���0y�U+;��M2[�r��LAͷ\���e�#��>T��a2|\�{�7��ә��ME�eiO���p��b�(�hx�Y762�Rgkt٠2e�RH���F6)��6�c��uZ�
����Z��}�<υa�(�Z�K �<���A�x���*�/;�*&�&��v��(��pڸY&�>���N0�x��l�g➭kq�_����L����(�E�X]z�߄Cu&��T��95�B<<�ڈ�~W���~�l*k��J�?f�-ź���!U| �G�NDxX��K��@}�"qw�C��"'�\��Rg�D��X/���<��I4�Q��z=�өW���R����i���C��T0{����'�Dh :�}| �l����_O�A�p�v�:8�xK�ny�]�@f�/�v�L�GLk�w-�2~�F;ҮR��X��K���j̒<��`����"0�Wj�q�x�|M��e�w,4@W	M*&�I�+g��u;�F��'�u�����E�iT�఼�k����p<�N���:
A" $��p1��\��b���q��h#,���7ꥦJA�7��Na�l����3a����J��_��P(��-�Z-X$z�}su���� �x[���J]
	EqP��BJ
7��_:�FQ<��p��d�E&X,7�bG�~9�P9�Z���6��2�[L\R3����2k�C�*;�)��ޝln�y>�gGy�(�Ǔ�i}��۷�e��0��%��Ã!/��� V_-�3ˉ�ul8s,�3U<:�v۶�2��Q���!�K4�$U��g����W[�0ޕ�y���T��F�Wo�*3o�6�i���<��^me`p�l���e[2�z�2Ԇ*��u�����=ކ�\��(�8 ����g��z^lñZ�j�kY(�D[�	��Dj.#�odbf� ����F�f�(a�vM�_&�1��I��B[�ݎ2Ó���0;cQ�eI��55�i��V�뿬���@�˾�9�����T�p�a�.�U�J��������)����չ�7ZNc��p�T0�AA��6ݺxPMZP��yu�����\�k�� �N\�4�ɖ�F�d u�?���4l)�����F\��z[|۩%f�����/T\��$"K�v:�!i��7��}<g��D���O��5Q]�nA��6�m�������j��7�G�=��'��Z�^�}��5.sp�LU���ژ��F1I��*�Kj:���:`"�����(�2��T%�����/?�<>wD���-�W����6yOMH��R������$�Cvv+f�{1>���GB,6��WSQ����f76�R�`7	���{�b{|�f��ֱ0���E�ҩ�`*��|����A6�e�;=�����53ݮ��t�jX`�a�/A��T,^���{���4^)r箲��ߞ����0Io��j�k��O�,��[~e��d�n��[� |�����\Y'(�d�[�u���z+vu������	�Y����KOZ�Ć��z}�_F���h��l!/gܻ�yk'mA�Z��������7Ʋ����O�S@b�J��b#��?���J-B�CV�>������_��oM�><��h��!i��}n7T-�7���w[t\ڀ$Hݙ
D&�i`�c�W%4�u�	!LQ�Uj�(MV3AV�S>U�D��Z�>��Ή)�gS��?vq^8�⣀�<7��a� ��{jL����Z�o<[�:ɘAm C=����pY$��	�ܸVe�V�J���|<�̑�*�y*��$�ȫ�� U�C¬9���/�BS�f��摯N�<�=��O��9T�P�Y2�h�-�c�7c���M��K��!|���Pʾ��,	��rr���o((l|8T��(��zdǈ%�0*��ns��4�
��U��J&|q��Uk�Z3���X�"�����(����}���cP&�+T���>��Y�4]sp1����3݋���P\G/���-����c����[|�"-/AC��-W��;q�|b�$ZD�@k>�es/]X�Z/�����4sM���L���6����O$�(Pd�և�2��V�$�q�Jq�޲��(% >R��1���=ݑΓ�=Ÿ ��Fo�{pL/�J�*7X>��Ql�&�	=~�Aa5o�rGޞ�|���R���-u��0�T�u��[�̩���lĚ�빩��K�8��h8J��"�5�������&~��uN�ΫQ̕9LDT�sE��f�."R�XWH��a2�+|sW`bN��.L�����_�郒�qX��B������̈́g���aȠY�'H� ��M��rnJLĄ�K��e��EL��22�dI�\�چ>���!��^~�E�d�hw�J�~�-�x�@>zj_Ƚ�N÷ y|�颖4����^��]r�0"殬�g��]vy�_���#�����j� �j�+������`� �Զam��&��!?�0�8��4�Ř�Rz�i�TO/��]�)�$\��f�;K��X�5�Ʊ2LSu���.�
�H��[0X&���.��iZ+cu�����kP�.fs����b}��1�X�|g�ѾNTD*�K�&��	|��>������b@���_Q���d@\���:Ez�36��&'򔼣�P+u�ʁ,�Ls����!��{���ƩI�Z�*�����XC�a�\� ~�:�t��}Z�pXl�}��V�O6���x���c����R��w�U_��������*�-H���q�����`7�i[M���,���\�QS��S�la�F)�����[���^�ؽ�v�U`�v��'����32S�_�x�E�ƔZ��qSU��Ҿ��>�>�����P"��?f.���u�'Y����cS�,L�p�"w��G�>��$o ��7����i���D|I:�zo�x�.�RrJ�T`-�wk,2���K���8�y���AS�=�'U`�J1�P���ga�ǣ�{�Z�u��N�����S%�)m�F	G�K���Wm>�#��.��lTM�s�to��ߥӷv�-���H_қ�4��F���,.�$T�/>l�"i�%��k<��ɠ���!�e�^���m��9�_OឬȾl��=�� ;J"�ݮ��J��b���j���;�3�0R�<�$Ae�?�mt8�Ȕ1��Z;1�.�x��G5��`a��l��w/�����_S܅�L�?�H^��A�uXBDʊB�=�S]N�a̚��er�*ޥ
p��9ěK����`��?&R�b��S��t T��K�3�M�X��� ��y6��i�f#����[����Bcj�I%䨓�3^�<sf�lCC^��a����I}~5ES*�]���)(��n�"�G[��;��,��:�=�1 �KZa��+�5��o��?7۴��S�FK- +\�u`�����~��a9��]\��i�R��<ůh?t?a�4@�N�7ggx���*�ʅ�M��ܻc�������#x���G�_w0}�6��8���0�U8y��s?�:
Y��6�p�,��M�iu�x��O��_�u�o��#�:G�TxAqC�7kz�e�>R�;�yk��#��l�T�ҟ{���	�$����C�)�
��^=�ך9em���7<��"�r-Y#>�%��H��0ʃ�!{z��s��YfA����7��VI�7%d@g���1dך3`%�����c�^��[��1��^-������D�����"�Ҿr�Z/�l�g����K#)p�S��7�x6�}/�2�J�zm3�0#`�Y��^D�d`!v8���=����^��jvӲ���~�=�S�8���%wd��ؕ�����}o�ck�m�$Ξ]��1-�+}T���>C����<Eқ�0�/]Am+��S��]@N�:f�����9������aۈ� Έ�����ϗ�e���NE�#"o�}�.v��߃NR�3��cw�
�X�����v��X΍(X��U�lO����o3�(�*Z<FO�HK�/�z���H��6j�P/&hN����y�(�V{�fc���˿p�%Y��c��o��v�H�"��M��p�� ���?o���[�S���Q��׈K�)�Mt���!v%p����F.ۗi�-�����hyOE����k���4]�4޿�̮}5 >n&F�O���͍l��F�4��_�����X?,q�Y�i��=,�>>e��u�Q�Ħڐ�3wT�m���6X@�7���e(�sMA�q�y23 ��B�-�E�����06�g5�d����i���~��m�U�ńc��G߶�p�Eh�!�*h��0'��/l�ٞ->N]�m�M��[�e�lTCP���h�>��N�s?|��9٧U�By�U\�2��խBrϩ�;���a��mهԜFVYhb���}?��+Y:��=z�W�Дz8�DB_���݁JxV�%�ٛ�MiK�bp߫>�m0�m�p	�P�T~5

�Eu��}a
Re@�Y�Y��2���Jgw75�hO\�Q� ���q��nnt_�`ZgB�?�׍#q)�*�50!# qʲ�D�#��t�RĒ���*�Y?'Km*���|b���cV
��[��H~A;�zBZ�&h����1�>�q��ψ	��Y��,f�v���IS���V���է߭Cv��c����LM	�`&�!x���D�em<i�2�E){K��2�v�ٌu)�՚2$��	�e�(�� �<ڳ)�Z�F,]K���y#yS?��x�ûM��.}i��������rw�G{�R��m��A'N����fm�m��(8I:$ݳ�h�1k5�L�z���<����PM8�̷_�u������Ό��$�K��p�Yϖ����*)�*�:G��ݞu��`�����M�1������O���<瘎�€K�.�rv�_���Qn���28Ɲ���`h��T�l��)jz�R�xF(�����dy� z�s�^>ף��B�j�V@�R�I��7���8�,�<]�A,�����'�2s\�Cr	8�9������3�P���1fsSv����jQ��	�̔�%yiL)��6��o�&���=/xj���|~�N��+�ޑ:رfŏX�1�K+��]�l�3L�?Y��y�!�%�#�{���[&[��Z�/h0��p8�r_L�@׃�bTdJ�ג �H����D�Wg9Pt�����E��H.:�H�N:�n�Ρ���k�GY	���q�e5��t�*@8Xfa䁘�Xͺ��,1��>��l���O�0��W	ܝD2�]�t|W� ���\�F��(�]����XdG$ow��<��|(���D�����ٽ�BP�D����ִ[�Í�O�U����C���>�������f�E�s����`��So��w�ك�.m8������A8��IF~gVs�Mnf��P]{�}�Pߵ�t���ݪ1�j5�˲XH�#nI���<��8zZu(.Qx\PU�Z�L�a�B��v�E�M����SH����t���Ú�ު��?����Lw�J[�g�@S����.�<�l��P&��0�z�f�@�m���	pZ䫶t6W��W�jv�i��Mj��ޖ�UEG��6��RCZ!�Y�Rޓ7}��z��&i@���܌v�Myeb�38r���lzp��
�%]�����n�R�J��N��7���UP��זhG��zD��}[,�t�)g����?�A,-��S�8�A�f��9Q��*Ж���[��#��{b,���Ι��U
�\�g��cV鵨�k�7=�s,�����Z�S.�o��:� $�5�i�	e����1,n�]�d����� y�A���gE�t�S;��:���O�����T>�<�U��T��E�h1#@��Qt��Xq�GN��{�~��z*�������k* ���hr4K��kW�ԥ � A2<"��BΥ�> Z�����S�jfb�,�U+q�|�W���?q�k�Sa���+r�Jm�_����x�{�|=��$'�֢^K�ηڸ�^Ai�,Z!�{Ҟx��tu�J���߂��b#��7�(R�4� �"m�>�g�}[yO����%����G0�b?9�(�ϖ����VF���B?f�P��7��x�MB�~G��	��G������b��W
0�C`�3��C,	�Т ��F�/��9r��h�"kg����7叏I�y�o�Yk؂�:6ۮ�Oj��a�\�t��p�]������<�af��B�z����u&�­�,�U��*`d�1]^�8�{	
q\\�]|		H<��{���g䇣x�r��F'T4a){J���4`�uy��j����v6�U�M�����4u�<�<�����"ȸ�SL��3K/]qq��T�p=\\�/���ki���;@U�6�^Pm�|�cQ��]����ktBih���6ؤ2�����^���v��@j�<5��K��V�4�2W>��H�Ӻ����~�)f�ĂH�ce����|k��=߲vQ��ǵa
g���,f�,.8M\44�{�A���mkԣ�hv�����s��,�w^O�(8+)�g�� �e���O]ŝ]?di��?�*>��2Q��C����EK ���ITr��_/r7�M���j�پK/�뫗�� q��� �#�D���	\��Gt��<ͥ�����G�%/M�|���d��<%u�A�q��5�K�OzY�u��I�-ŨZ��rv�LO([�&im>2y�qq�{%����r�QUN�|�]���R���mf��zg,��䗝����I-Z���x�%�V�����j����ɡ�۽��C�v�2F�m��Y�>�$'�P.Y��;���8J U�"ɽ)"�~38�_!�]��n^@�߻�a"�,��sG�w:�nU{�UTS��(?]�O�]�q���h�3�7��.�H+���ʝCX"i�}3�˗'���@Z�>E�ՙ�>şQE���׎R�*Q�k5+�i�;`������z?�����=9�l��/��G�7�'{��ړJ�:�U�6K���b[�R`EPh�;X�3к>o�[��^�>i J����q7X �N��l;����D���	g
Z��a��g��'��u>�����&;a��(~6E�ޏ��C���cx�E��(�M�_r��T���zқ�'[�=��`���u,���	Q��4)=c:��	-�N�πo��H���4�N�
ϕ����}��]�u�����N
@����B�p�g�g�T-S�0W�Ӱ��E���ߣ��@J�Y4��ʜf���ԷmO�j���0����zV~�]V�o�zE��]i�/�I�R^�y�靋)�>�_���טD���PI~nE�e��gh���b�N�t
�q�'�8��&$��ϣ�����|��US��O�����H�A�rZ��>p�rƔ�:���D�}���n ���*ۣ6����S2����f���I��:feѕ4�_-|"s�.���Sth �[��@t �e�t'�[?A���Q��f��x04�:o���u�Q�x���Y^��2���N�g�q�a'�$ T]aj3���(9��v�Or�0r����k�*���Zc���}̄&��a�4C��|b^/�Jv����V���e��<�Xrqim'��sؘa���A&:��f]]CУ8�Γݚ�\H�B�˘hؒƈ�;�dy+��]�fB@�6wu�����ŭ���U�n��#�\#%��%�]�*;�Aq]+Sɪ������� B�Nw�؛v<OON�o�hZ��e�nu#�N�@<�L���!��a�
T1���1�@"��(7RѢ�fdA���ɦQ ��e�EtUn������x�c�;�R1C��Fy�,�<��D����A3c��j��b���ƷI��@5�ҹ�����VVwS���7�ӓnbw�#!���i�+���Mi��]vu��I�x@|���;wQC��;'�5��v���L받�&��L&̫.�r������r{W2��&�tZ����4G�1��Ǎ����pDڇ=��w�������%{Mߖc5P�(L�}�"��\ͥ?��j%Tm㏔>��3Jz���(E���o؟����$�?ڭ317��"c�9�Q�?�LX6֋m������E���cu�'��"VPj6�����3�gڑc*�;�Ϥ�_�����d�;��aC�ϛ��5��y����떎Q�V�BO�	Z��R�Jta�:;��K�@�Itzd?�>�ǚ��U��}E1v#z���V�-E��_8��Оp{��^7�G��b�p�e���`���C�k�n?�cK�n:�E����ZD�oC��ӉX�^�����s�@�$����g��c�5]-��;�U}+�JǙ
�L��EClT��G��P:fV�	za�sh��
�;j(���ѣBT��J+خ�n���+j��-�y��4y�3J��W��^��7��O��m};^ �l#��r;��C�׮�R��_��ɧ��U��s36�4	�p�cE\]��3����,��3�u��E{6?ǖF�Ǆ���i X��37��fk�;�QV;-{�
�~��*�3u�S�uEm�|wacfR?W��\u��wd�	G1��4�hOP�%V����\pu|6
P���ޕ�G���WD�-�;5�����_�d�Q(��0u��n�O���3�̵'�âa��55�����>I�$�?I�>���?�n���k��c\����fyʈ:&8	����	�C9���M-mQe�Y&���$�����L�I�RQ���+�i����y��6�畽evSN�ǝ;�.��\�-���ac��|�J�:�6	�F	��=*I/BC��8����ɨ e�zUy�*��k^]~#�|�ºpԪ雗K!��뷋��!�Kz�D��>`���FƴP7�ЧR$���=��	;$	 ���l�w}	t�m����@�|� �o��S�����׽����܈�BE���c�a�{6 mDAPD1�rQ�Ydה���a���)2^@�A!q'�cS���
/{�Oi��ܦ��9�U
y
�]7����V�J#�P�Så}�x&i&�*R���?�������������4u���)�Kh2��uU�jMͪ��o���ې(������T´0Q�b���\��?��#\4�����Bp� <Q��K���_>J�6�p�!���(���~=@��}�O���G5��_{���e��ό��f���faH��8�.�bn. ����d� �T�����<9�0��э_� ��2�8%M?���PPrJ&�e��ͪk�N^mь0P�~u�g@*�ܶ'�+�����,]��c	��3E�^����/���>ն\����V�b�$��s�h��2����������@��V���;p���g¥�%9�m�	r?�T0{9���^���>I<|���)�9^|�6�G��p%v2Ǖ������O'�j��E�I��|�Ұ#��ا�|6�YS�0�S�F�7�}�d� �u{��F�]��A���7qlP&ɶ}�v��6au��2��� 	jv�dp��A�T���]��]I�׭�Wl�g�urW��%OL��u��ID�-	��ŀ�]6ZH�x�\@�F���ռ>{��M��<��;�2��Z*�8�b1���^�4�VS�`aS����DT��0)�
����[�&�6!	q~�<�������K���ql60tt�wfUg��.I�<S6��Z @�G�ъa�(�nV�#�+��^�j�b�4Q�u!�[�ӗU0��I��[��z�5�%yK��x=T�M���NJ9������$�G�.s�P�jN�\*���sb%�wp�����?�ɀ0�r��:4���.�����g��@c�JNm6'0vp�]�C���}(��˽�$x�������8������Ê�6��(���V���F%>ԧ���Z��i@����?�����
)�XXKY]��讈SB� Z�̧�#���̀a��~F�KB�R�4�_Y��J�ȋ�}6q�C/���{j8�����a�!\��Xd֢�,اp���e�G�=���=)��O�c�t�&K���0��r��
�^
���\���$鋼Ը#��TP���$=5Z�1�'��ل��`R\����������Y��1���t=��2�j5��oG-K����);��uNvD�H8�N��A*t��?� ˫o?�X����v�N`ռ��*4����د̜���*Q�����UB�R��6L�}�iܼI�P�����{��ɕ]���Q��n�����P�R���ޭ��|�T�^�v��{�.��D�׶ӫ��շ��n��醯��0�������2����(��F�fV����l �!�}�xٕ����1�&�=\�s�@�ʉ�c�u{e�����ٶ/&s2״1�����[�@OZ��yE�=��^��Ō�2��A��Kvf��im�9��hf� hq�U�搡��|��� ����zR�����w+,N��\2�sk��F4\��ҷ�4j���g(���s���:��}
�װ$m)Xi��<u>��)6�?��f@p��sim}a� }������m�F`-��ԛ���cy[����O���m��H�$�5}h�J��\��y8��W<wm�ѩ���^�(A:���i��SQH�d�eǀ�0�־�"�!�M�x��̟L�OOB���������ngF�ή\lYkN��̾���GK�i���,�'�F*�3=p�y����݌ O)>b�챁f$5����-u ak�i�����+�3��u��	<���Ash�;�9��Z|)�̺�L�:���O�s'N�w1�mO����f�� �������s�̫���
���$`��Gtn�/e,��HI�n�M5\c������Y�i�8�H2����v��^���"�s@O�(��V��-@L�H��M�.��Ƚ:� �B)��֕�u�z�4/A$��1ν�\X/��U��U	��D:�/�Sư��s`g���b(n	���Gq:����	?̗�p@��lX�5����B�� -���#t��۴�H��l.���,���Q�jlH��o6>2�UQ�虍cd���_�~��?�"o���G�sUn��w�;p��O0h	�ȝ� ܆;�H�"�H�t�����o�4,[���B@�%cH\]�u�Ð_�|/��B�ѬQ}jg���G)&�4o?�&oc�o�h��C9�`����ݡ���^��������/���{�X���iRI��Cé�@a�6D]h�	�
7{����K|�T�c�٘���3h�d+���N��'QxS�K�0�4c9(��L���_�Ϋ���3N�>(g����gAuj�i���|/��Fkc����7��S�y �E%����9���ԧ�^�C�[$�آTac33�7)F��ɱ%�]�u��ȋ����D�{Z"���P��5+��I�E�s\��l��3�4`��{"�`�
6 h9��&S H�k���ə�?�Ǐ�g)��(\�]�Ђ��ai���f��_��!п���n�2�;����cq5��Y��a�>�%��o�J��p|ܳ;�&�k} ��5h?�/}���V��}К����L��Eepqf�"y 9�c�7ף�f�4����*o�G!ކ:�G���g�*`8��pn��J�!v��^�%a��ti�Md�����(�6'�p'�c}��SJ���./��ʙP�^����.�/2g=u��U�˖��3=�����@��?Ž���FN�L�쟧 I�I�^>_��^z�(��V�HE��tE����?G����Rv�&�XB��F�������%�3Ƕ���oBc�9&����f�����yܒ�E�J|����s��Ϥ}�BS���%Ӵ�����3�p�5��x����l�e�W��^�[���Јn���ڴ׌[je�i�/uN�+[�� �v��v�6j$\b��w����z�I~�ni���c$������ t��_�H҇4����N�T!R|W@+cC7�r
������L�|:X˷���OAވ�^>r'�f��)���7�T��~E���`i7���ő�����8����D6�TϢ!��+�A�ԚJ�[Crz��_]X��V�P�4��m��1�2����{W�
��r+3~7ZA����C�ܣd[Ǆ?�,g��`��\"R�����d	�C*�4`E��οЇONK����	_$N�����k\���0��u��^���hU8P��wBs��M2��l�r	Ͼ��� ��{|�݁O��s��SW���֧����<F��Q1ڄ�#	r�p�7��^�w>���͙]���a���?p�X���wӲu.(���l�j��s�����3[�0]Eh�@f���r�"��g@��^S�í9�!�qWoyf>T�D1Zm�fOM(��M�G��MIt�#�y�_���y=���v��POэH]MWE���Q�
��V���0��|b�ˏ��O��"��aCm���1���>o�w(�E����vxGȈ�q�+F`э�o-�'V�k�ho�/J �[��qy������EV�ݛ�� -�X+���&��T���\V�~Ur߯Pe�pX��1��?Ao2���[���t�0ry������T�>�v�(�#a�j[��J*,S=�0n�J�ғ�mc���SY�8s�C���ΒkJ&�������DA�2! ,{�`oqMU�p0�p+ ��$��@���Q��4�T=&����
ҫ�ڊ\�+�(*�7�fi.������Pa���x�#�b2^l� 6|�@-��)b~@F�"�=TH�N���ȋ(��B�]l_�fU�Oμ��� �<U(�;�q�oY�ܔl#h�
G�
��
l���;5X�P����B{������}���D�V7��}*�߉�"��s�d�&��ԶuMΠ�5��_VV.�����zq��vv����U!�x�~���['���5��0 �yݑ���ԭ�/��\Q�.&u�I*��L�,f�:�t:�C��hs`;ޮnb�p�˦G�Id&�F"uX��h�|.�kL�-�V�	|VO�,�C-���_
2�𯜜G�D�<��_��K��޸fy�iW��T�sc}L���&	N����@1r�EӹAou(%c]�*�Y� 9b�;:4~l�H.�R��,Z�Yv���n�HE��g39b�hƺ�<D��=�θ̿�i�:��n?����"�j" T�G���T:q�<�k�k��$�U=%�vV���,�:�)q?�_{�7���L�5����JnPL����239���K>�DJ�!�1��b�\!�r߆
�[Q�J̑ϔ�$�%����y�[v�������N���6�0A�J���X��
�%^^<�IiIY�x�4��%�+Z�6��0�+1]eބ��/Giuо�U W���s� �w���/���5�n�~�+�?H��Vz�����=LI'7A+�9Z�*S�S����نJ�s�k6"z�~�5BP��5Ł\�j����fDѠ �4U���U��y�_^���	�����_w
ӿ��R�G����w���I>!��XR�0J�<I	�dPz\�����zэ!sK�Z/(��� 4D��
��������-��S=��`{i6��M�YL�P��)Y��W���ܿ��l�;�0Q(��O��i�Q��3y#g�m-{9s�G|Ă#�S:�1}K�]���8I�-��P�V;���r7�:\�*�5{"jű�T�۬P�54�F)�v�}ۙk�G����E+Gy�����gK����E����q�:ݪ�_�s�R��1U_@��%0�*�%��*|"��{�Jp��B7�X����Z�psRo�rX/�������&^۵�U�DM�f�#~8W8�j�Pv�6��*�b,KG��/���L��y/����,ʝ9.���v�
�1Q����|��:B��j�b��+���~�4��W���N�� $5�n�+I���:��3q˂��?���Zl��E��"g�pǽD�h�1�X���}���X�,��+F�Y���⪡�u�,��@5�m�����K��<�vgH
�;V� �W�`�G8��sh��ù)Ɓ c
'~�S��0�E>��OPIIV�-2"B���j$��qͫ܌C���rw�vg�؁KhS��\��� �bS�`@&9`��6��4�3�7��-5cbzʾ������P��E���@�3�*?��cn�g+�ڷ�`:�4 Ya�C�pXSHQ�Y��kC��d=s��\F ����,SMt9���g�86D�i;��Iy�?�ⰽ>vQ��^�8ӕ�'�����Y��KV<�����\�?8ca�0|_�����.��Zssx�0J96w�	�ֺ(���f�M����N��93�')���{=@�s��Bp逸>As��2�����o(ex��@�Rnɻt�=���h��>��brd�d��;oN��`r,���aAt��s<_�mV�2�"M�b�PEx&�F���2�L7K�	��ι@���ܩr (��#�������P�JJ��`��3�t�h��9O}�M�b:]����������}/;e��wC�2Г3M�B�q�������oV�ls��
>#[dsr��
�:���]��14��D�@���*dt\��� p�l�	�g���1�J�Hy����9OЀ��}̏U"�fE'���]S���.GBYx���JITF�z��S�R���	4�+/$aOv�����"�f|�j���2����j�O^�V/ �[�<c�]m��E��J�ҧ�vO����z�y-�F�g��>�GG�k�����}5�qZ�j�=�c����
��u��|l�@Hcg���T�x�Y�p2Xȓdn�1#�k�lfh�:��1��;Ż�p Z�y��q[g�@-v��1O	=#\���7xr�4��qN���p�w+�66%u`s���esel���?R�����;a)=_ګ�i>��WMR9���Q@8�O��i�:���)a��k?q�[��H���~x��pX��Q��}j$����D1j�H`k�X;/��G�I�RZM�tg��ҍP&��֔�C�cj-�8t4�+�F��VzTٓ�Z�H?��	�5O~Z��#U�N p�}��1=qm0���}�����i=����%!����Q@w	��<^�W�2����\Ѓc�+HM?X��Ό���݆�O��ȚڮQ��a�Z3���? ��uaP�����Q�iG�Cs{bA(@��=��(�`N���c��@�(�<mR-�r�1b%�Da���&�{F�2�ű͋��
����Ҫ��� ��M~R�UޔZ�����Jw`)�����J���g�=������Ƞ~3ȸ�tx�F�rt���KB�2x�M��1�/;��$^�&��ok,���kP�0��2��gwg�!��T���:��l�����\��c��K����7m�Y+��8���q����uy0�Y��\�1���q4��*�f�3�$�߷G�]��$+!pS�}���IxHzܖ�1�������6���{�ɀ�z���ځ1↹�Y�T�R�Q�Ǯ��=��Z��.=������~Z�/ց�x�W��L9�l@�	wA<m�D>Y�W� �Q�� xT/�3�%�~U���+����&�9<����� ��)y8R���$�m��֚�x+zE(�d�������nF}�!�z��>7�[K(��pdRq�p0]󔙩:W$���z�������֍�]W�n�{<ǧ�)�z���/�c�Ktv�V5�VE�_2�?V6	��;E�<�gԖ����z�5��]�3��q_*�A_��ɾP��	�K�1t'�����XZi�U�h�0xC:���%�W8"̢�)Y�K����	v]�mOk���t���ɿjh����[w�����{�&����W�1M8��`4�A���Y6���b:��aB-_
�:E�#�q?i)�v��*>xk�0ج�q	y{���"�L�.}󬻣�2F��s�����'</�}J�J��O���!^�#>�o�YR�؋p���j,4ʒ8���L9wޑ��f�SG����X,.�#������&}�x^/�ueW���&�#������i}m�j���tj=��CPO	"�O��;���y,Pb������qȭ&!S�x�/2�@>�O�9A�>�-����!]t靚I��&-���YbZZ�n�+F����S�4���\����r��6N?���~G<-A�DR:�6��׎Qr����r3U&�&�-N�u�Qb�d$޴�Sa�`nb�-�3k����>�y�o���hp k�Q�vց^p��祮R��!(Ch���Ms��bT��W=
x|)�\xs�}ARy.�Q�� yAN3"������=M�@P;o�{žY��.����e�!F����3��f'���<$�By� E�I���n���Ur��u@����i�8��A*�=G](�����8\�o��H�ű���<!�ax��,/]��r��Ѿ��A�^�V��������8ы��mNzC���8���6)�A+�%�,���XnB��/W��<�P�4q�}����+:s1�͟@������������s���T��X�]��x�r��	�-�{,J��i����`b@U;���������&��d��'p	/u*���E�ң��E����!�ǘ����y�D�>� ���ѩ���m
&�h'D�^�S#�A|�}H�i\�5�14��\Xᒪ_*�Q��҆T}$mS�Z8����c�$��h����%>�Ͻ��;U�Hj;TKe�;���_k�gcȼN^Z���Js�xnm��yU,A���k��XQBn���%�MB幠!�d��D�� �N�	Ru\
+�M��� v������9��DX���ѯ1���������چ;;z��R�aҬ�ln�H�)�=N�$��;����W�./�����-�F�;���+��7��0�on��r�U��{i��� �=�q?d�UhvCM�1��2�Kuv�t�������'���m6���C��}�SGNt>6��AroT^�NMAc�+�[�� �� ��6W�(�K�NV31�[ߓ���{�?��#�?����l4�=�fīG��B>�V��c�,h>/���t/�8�h���4OhV�����XD���Z��x�gD8-�����H���C.���c���*�vv��tI'a��#���u�M2��]�\7��<eD]�g����K��W[ԟք�4�<�d.�9�|h��	Vq��A�b������Z��%S9��]xy�!�}6�/�u������ӎ��-(���Q�`����w�ԩ��jP��@����b���t�*V���Ҏ4���3�^��H�7��uv�߰{&�'3�P�/ȳN��u(]&H;�"y�6l�����hm�T8�x���`��Tgi.�u�{ȿ�Ά�6V�M��*
��,,c����!�7�|�&=p��&�3����T��B�%��U�]�A�)u	w�����_�������EZ?�U˶���|)��u�A�b-Oq��*wϧ������0\�W�ϐP
-ڭjd�z�wB�����#�SG$j�W�:)d��˧]}&+�F���/g�ʦ�=���ܚ�t˺����S2zxM�(�=w;���.=��Z{: m�/��9+4\�� ��)�a/����/���z�$���Ɋu�_�4t�. �w��yD�����
��u����wtiK�&	ʹ�n�r�~x+���
��GH.�M���jIm +'�dT7F*�.�d�.S(Z�Z�E f7&�B�c����ޥƪ�dvdNA9%<`2�0�����OC���|_���j�ƙ�Wp��s�q�+�)��������/x�z[̀���nx]=���X`n2��h 9]���)?R�a��ww�V���;�u���dh0�y���_��Ǡ�@��#ܢ��y���B���WHp�����F�ή&�W"�� giF�4%ǰ$p@"1�|-�� ����h	~���\7#�J����f���V�m(&�"o��f��u�������nȘn�m��nk]2��t�������NܥdIJ(�[�L��K�y<`Qb�{&i)�z O٬�!"	|_�Qf2	����|+K|u��&~���9�����W��$l~����Mf�W���"K&�h��9��^s��3m�B<ҘB�z�K*)�B��m�G��K'�\��,�7�A��|B��ұ3. ������c��U��jɂ�C'?��)���;n~n���e<Ne�?
c<��v�yP t��0j��������P�[��68��{d�L 4��v�{�(��if��.y_ d���ŷO-	��(�e�ү<�ؒ��G��	ch2���llZ����]������m	ͪu>��X���xi����*��Z|����{�(5<��\��"����Ȭ�P"�W�	kػ�5��1x!�H�ɭ����j�+/]�p��&GW�ؚ�ڳ��4g
����~�.A`�_��3��S�L5�1���A��6(������x�1!ue�S�ּ.	`?]l����wҲ>jF`�����b�T�Bj®��*`��%�$�(��V����F��q�F}QFH@Xav�^9���P�T�G�
qj��lT�!���iWA�J�$���&��������e��y~����S��,ք_�����[���_ �*?N��j�ǋ5�����gK��ƞM�;��Ȑ7�sj�Jy��1����E�>�wq�ǳ�$IT�[�U蹴� ��wfܮ~j��CN;d����z�r©V>>=���ú@K{^���K����\��KtU��|����L�ŗ7d�7�J����m��ylt�v����ߞ\�^h����ز����o��Dd.�PD���(B�/{�,H��F{�Kɨb˳����6՝��P5�����C�H�^}���
�d<�*��9b����y_Gӷ|?:B�rkjX!t
��r�T�� ��wI�NR��5ڜVN��J�k���� %��B�{1��3w����b�c⋣qeJ|�5È�\*�k0F/J��t3)$����ZfDQ��ddVL61N.釹E0l�	Ғ�|c�I>���і�j���?�f�d�%E �w(�Kf��K�g��O+Fj��Q�1�/�鰰 �dBi��ⴐ��k>��a=�2�;����&W^C��i���Mg0ĵJWf&կ�g8i��u�)b�Z�1�y�v��h"�A��_[Ͼ����l�=L͸���,f5�^�;��� �o���2��*4�]��?±���pFj��8]Ƨq�l�钪�E�����@}��TD���C��*Џ��-�֑�l7�Y��$���U�gð;��t��K��T0�w������p�V�9Bݰ�2R`�_�:~M,����ޣ�
p��Y	;(�14�j�x�k/��!R�9���T�լ�C��,5V���Y�H�7
A4�������vji��}4.Q�����OS.���~P�}V��;�Pj�ǰɲzVj�!�@Q����l�`"��D�q�T����*"w�q�6 �-B��䮘�B��0�����RG�"���k���J���߸v�*ɏ
f�y�!	&�AJ���Ĭ�#P�d[�M;�0�TC��z5���n����˪~,�j����$V��t�5�I���m�x{n�YQ��a_?T����
�&G��t�TU��x	3C=&��U��d�u|�9�H��_�U-(�l���Z���@�u�]�5������t�}}�K�1:�A�(kǰz��Caf�#KI��*�!	���R*} �����*b!hʩ��Ħ�5�� ZZ�&T�ڡ�݆�˪1�4nI��ʕܚό��60�*����%�NaN�͓j��xD[�Fݦ~(�\�E�h�W�>9<Z���W���*t+�����{���l��x\l�=D�s�錃��Uԇ;�EgGKQ=i�k]5WK��K�%Q���c�W��M�j5m��i᯶>���Ȭ�N����R�*dsX���zM4����'�<�.�/2���W��TzC8����P��į�:����ޱ)w=�kܺl;�,�&?�+�v䌪�;��,XU����mM *	�R�6�!�5�#&}1�̀������_��Aa^�Px��,t����IzU�|�0g$ҡ�?��ڷ�R����-fN7v5`~0_h��d����r�W��v�w��y�G��c�8������s>�
}8{N�����b�j9�p�������搻���Z����_*�A�M;<�\Ĩ��P��O�-3��]��=*����~T5>l�gp�Mӽ�Lػ�ˌ��wJ�<�Kϯ��V��/﫷9ὣw�(b~6�[tȫPj]($�'�֠��&�[�~��Vfm's7����&O����]�q����$�4	�u��3��/'}W�Go��%�Z���ǌ���n���ΚZ�8�7�����rVXeo/�R�Miό\�5=��K�旽�O0�=Q�'^�ĸ�zY�����J����vX�h��lb~C!���C����̧�D��Ȩa�e�����Tyь��]*���9)	8`�o��is��.�g���Q$:���7�F)#�W���"�� M�Ӝ�-��/�/R����D3>�}��"�ꬁ_t#�=S9�g�5�������������jq��N�4�fna %��=�G7z0BzL�c�:�+�}��6�/b5U�o���
�լ��L�;�d�*�r�C�kĐU8����b��\�Sqۑ����^0���EJ0~���.3��sp�N�n���n�wC'��jhhO��H�(�`{�7����\���IOs_� ���N2�rZw�|<��ʣ��G��4֒A�����g�N\KL�@��^�R��DG����&<떔��V��9̒5Y-(M'��/�n������	h�0J�=L)5�	�)S���O���Z+�o�HT[V��o�����+{�jP��*���2inUټ�q+��`t6��}p��y�:-�����R��-Lb�I:���6��i��U�EjEate�}��5�wv���2Gu`axӵ|�69�Z���EvU���R<�%#h��3ge����� ��������hxc��6���.? w�Hd����*�tA�\��Dy
�?NLN,	� �"�R���y�#���j3�#���ʌ%��{n,k�w��쯽7N*Th]�"$.S��	"H���sz�;(��g�5���<���,�K�E���j�OM8��$vi�2�Ŕo`� �!:λ�@��� ���f�8��N����u��B�\�.��S�y-�#5D��x��Ɠj8�ޛ4X���xK���O�]z w�R�3E�G�?V*A���j 4u�6_�B�w�%O�R�G�V�z� �<�	�r+M�N���~1d��os�F�^|��?N��w�r�����E�Q��©�<n�ӥ�� kE��N��3���A�U�-���f�W.�Ͳ����:N��m3h.rj"�[��yj'DĈ˕�C��F����I��ę	�z��n����ꠍ�-����r�����V�m��D�	����O�
3�L�?W�"�����EG\u�[kX�������������+�{�����f�c��_.|>/6�l���?���?|���G[����f��1 �ؑd�� L���%{>9H��Z�C��4cLM�*������lD[�%PiO*Z�!�7im�l
�(����>
E�<�=��,!5v�$�љ(;�/����s��B�*��!��Cr�1+�t�a-e.�X�e_oN	ftU��@�I�KA-O0}U�"�#yxv5�W�~ޗ;������l��P���Q�����}����<�b�;Ȅqx
M×��RӸ�6�3�Ι�����H����X��^��To/�]�Vu��M���}�]�{}���4�%��w"�������X�Bnçu�y�?+�fR:m��"v�c'�Rx>�X�g�橤1*�r5[���lv����}�_�4'��}�����F����i��%dh�Om������
��\��o���8���J��La,���'�)�H��ԫ:�\خZ|�a��m����~�e��Vv�U�@�Y�P��K�hJ�gRb��@P��=�$6��O��$�^0���G��̒�L*L�$����͕F������Uy4������jI����*���l��{f�,$����@��D���������0�"%\X�~�H'(�POz����Ë�L�#��j�B6�DO�hıh需΀�>Y�����#Ћ�%�/���Za��3�y�-�x��)����h�%��ᝣ�{�h�с�hҏ����G�~kL"����¬.�
�,~�l�����0Bκ��s���Ũ�*�;�����NM�g�f�`u-ky�|�1�}{�¬�J
�Ft�
yi|��i!NC����)�[���E{n�T�Y
�~�@��	d�Mc���!��۵�}�	M�xS�4��&$�G2���:�[!9�������t]�KF#�u"SG(ZL���4��b��E��i	q��n����~#l�ԣXx�b�o��r_=���Tq�QT�/�����^�r$ٌt�h��9ʋ���=�5�W��N�
;<T�#d)(�ѕa5�Pow��Ar�؏`��;ۄ��lF�~�Yz)�bߥLրV҆����ك bbş������sfv/���f��D?RQ$fb�z|�SdU��^��|��1��(
1{��a���+F�~��)K�����x�y��Z�n�z����3\��r޴J��}�I�BG�-���@(��ۥ�礕��Y����W$'�l�˖��4g��k�iE�No��P{�P�8�Yh��%'\oA���&�]�Yb�G'�U)X������O�o/x徣L�2�V�`�����5����q��9��f�	$�t�#�UF<Bz%��f�޲Lݻ��B֥������r��9�/�=��;���jY�z[�U��	�Ԏ�h�>�Y�>?��+X�D��5.*�~7�A����T���~/Jv��>�8��M]6�-�t.�&��rK����/笐���f��T:f����F��y�j2���Q�/@�E3Mm�����=]n?{C@uƚ��WH�@�e������ �JP�T�^����W�-���:�;�#���[�vG�uQ�E谏}Z~�J���#���P��p�n�lk���1ͧ�Q��"s�ƌ�~�e�(��L�ck��T��1�s� ء|Q��6M�������g�n�AV�2���-��<w6���0P�Wڗ�_r_�.R�.��%|-�U)��h�Kn��{?���āK:��I�����9I��z=�Ч>�n�c%h��@W*`8n�D�X�^�h(��'��g���e�4�r����1N�c���L&'���OI�Gw�+�,���5RYݎ��vK��+y�N���1 ��s�Z����y�M�\��0936.s�N����=49y-/{� ?��D��鮝~�ω���qH�iҟ��/���l)�^4�� �O����{��h*5����مg#F�6>�CW6�����K��P�D 9Octr_��*$!�s�H8�� V9��B��7~*�,e|���u��j�7������X�)��i1��PG����"*�o'�`$��7#�ѯrW�K��-�z1�B����V��Y�����+e'N^Y�)C�� �E?�Z�濬Gs����2��,�0��"dׅR4�끺�F<bf�K�zZ2͔�E���2�jJ��W �]`������W�ֹf���_�N�}�G�f�o!�	��~KW� 6�ޡ���%��*�	�V5�@���rK�,��EA1��*�X�w�-����ܮA	����H��AX�������Ug���d�
���\?<O��S�k�&0T���J��$#)e^�t��+p���kΰoA�v`8cj����S�b9ݼz��V��^�>$��I�n�G]�[���P�{t��{�/��/�3��Ո�w\f��sF���"�Z�篰X>#�J�PI5� FK:���o�E��'�Qe�pE\����ލ�9p�B�S[G�6!�q��{о�&(
L�r�|��Z��8�G|�%�4EF�]�X(�k'A}}~�fc6{_R;��LMj�����F�@i�x�%�v�^��d3�z�݌��8�rQ������\l� P~1�0l���F#M�3��r4�h�/�̈́X2�X
qo�ڞ9Ye:�]9̴1��Fκ+�g��sI&Ȏsw����K�s���dY���¦onNi[����h��6)��2��6z�bgW��e�F�k:�5��D��@$�+�2�[�/fk�\�H��ܾ�!6������F���Fӝ��gDD6��l������s��{֎�
�*Au.�vb:Fx�'HN뉩��c6*����v��P�����ݶ��H��Ƿ_b�����Yƙ�x	���_UIL%���MHj[X�Yp�d�wT��(T��֦�ilJ�\c`��aa0/�{�眆߽��CB2��v�<.K]�� ��te���,xUM����@�{��L6[�0w��t_`����a����dp���0G�F�������#M���k�0�H �;�:��:_�qd�?��v�P]�ٳ��\?	���*4<�q�}���q��v�"M�dH�6@b�?��>'Dv����@��# �DY�5XU��*����'���#$��.��r���&�.ːU�z�i�TW�ՠ��[�U��tg��N���J����CZ"+��/�!a��*�ws��&rSN^Ӱ`<1���׆>�sL���Q�̿�J�\�Y���������ٰ�Cr���Z��D`i{΂k�.9�(7��Qah��\�MbB��X� �f�|�����]~��G�%�K
_�m���Ĕ�n4cdOlV�������f��_�#��.U����k����5pj�'BZ ���[������%S*��c��N�+H���r�.�D<�?�ڽ�#�17'L���R���@�2X���"_�4�v8��T�����Ů�(�70#��I�!bj��A)�0O��BW
��
�1���Y���5d�P,
��>eQe����>�%��Ț�S�O?��ᔾcy��5���d�+�*����(�%���2�Iΐ%U�崄X�L[�G�$iőɓ�v�Q�������Ŕ��`f��7
��.}'hi�v���.�ŷPwQЕ�$��jv'y�6��*+���7G�)˟|��p"1�L$r��rȺ������G�c�o�lIu3{zx ��,�K�<1��<NXlC���MF�}�#o�o��=0.^�v8/L��ը�E��-�n�dh��j3�a�"m�?Y�B�\��X[�[^U,L��.�_8�/"�����44޴&`B�gL�{�$�h�&�ۈ�m������c��[z�N� c ��>��a�32�7���/�[&'�U���R���k}����0�\sǳLy��E`G	��_5_��亇���α	:�L�E�@�8 ���x��NZw�w�)��
*1ʸz5M�+��s��uvO`l7����㍒���s��)sv���������М�M�;�f�KE��b�h��@��Ff��rr���y���ޙ�9�Z�.;�����<< S)J�i���b�N�uS�zGx~�r��1�yf��"L�EL�

X�.o� o�%�gx���C�V[qu|���z��W�ύ9۲ `�v���v~�h��i��Qʩ#ug��d���(��'B��H�
��r���QP��=�c�:u�P\NTЭ���Z�ay}�j*�$Ł��1�G����b����R|�d���fZ��t$���2��.�C�R��H���!S��7�דQ_,����Ǟ3���d�6��qa�,P�C.	{�\�f���'wc��6PQP�$�5D�5�������y^ �.��$�о�U{7T�!#K�o�!!5��٤`<|��V0�d$��SrT�r��><�(nފ�[i�����f �E��'�����������*���i��lNY�<0jCY�0�������[��s���|�7�X��&�y�Λ�������lLdiY{��
OVFώ�(n髚�Q���=1nh��)��]n�{�G72*���^HV�r��P�Kd�^��Hq?��%����$�X;�o>x,���>�����/��	�(
>��	��C�$˪X�9�(P�qK&͡�A��ܥ>��>&']���~_���7��V�
��5D�|3=ey�?o��MU'���|�����Z/� ��=�+���8�s�l�Z��9�?�f=�h�*��a�G�k�uǱ4�E��S���g��غMh�?)�U�� ��Ka�m�I_��f����~�A��+˜��1ލ��̪2�yU�D�lU�:�V&�bQ9��F��[���8��l���{��^��� ����H��T�=��UJ��W��S%�\��.����6ue�\�6c�W]�<�u�@V�����KD�������r��������d6�F*��.����϶���A�[�����G&�N3���|�E�IȮ��=ɗ�cL*;4��؅6��?ą�y��˲Y�ELf64��t��x/�_/w�U����`Vݼ���b��3$,5�0���,��]�Iʤ��@4e[��G���ya{��3Q|�����{"��8U�IȤ_�ޠ�/-��;�DW^y��0v�h���st�(YI�̪�Jy!�v"����<M#f��C��KD�*e�8��q�y�u:�f���_�B�	�2���.��L��t�y�Ҹ�Jb���rY���+i<Y�6���Yu�"m8Z��]�ծ<
?9����Yb���zx�UaK��#j��rh3yRcQ�i��E�T~(�۠�k�Ha�������8�������xcЯv�iچ�K�Dt�.VEm�Hq+��Ӵ����e�����M#׶�}O��d og���o��E��;���kJ,X�m�����c�7s�B��/��zW����jA�:��OFvW=�S�Y!�Ѥ>dY�Щ�w|�rvUK�,��u����*���j���)Eh�t�!̓]h�������v�s�Fs�����ׁ �܍���+Ӆ뮥u��J�K��Y�t�O��UY2��g�*6��
+�\��Χ7����d+�^�g��[�H|�7�(K���K�n��5�����̞���)"k���Sq8O&Lz31���N���YG���|?���0��<Y����;��F����,�D�V-�`T�y�ލ	F�f���Ļ���bʤ�O�V'��R{�bq���X�-��͟�m�׌�8n��z�w@��F�F:�r��d�i��N�<ۨj[�eO�o��{-��g"� �g!ꁝ!���6!�*�� ]%��@i�K���;G�T�V'e~�G��u"TWs����UQR�����R��#�jI�=�ݧS���x�	�9M;,sPl"v�]x���n��]R�L�Z�L���Blc�[5��@���k�v
�Z`��Er�\�h%��p�ˇ_��hv����J���:iv/׫}d�ڨ�2�����@����u��=nK�i��&4�������8���+��:ޗ̈#;1��S�E�c{��Zv�udJ���l��];���8=��#zO��v��.��I����9����A��W�����Bk]�s����vt`B����%m���j��Sm	(중0������aj��~�p�p/��r��'m������t0xs8#�N����A �G��������%�{SQ�+Au�o|I�R2N�)�F����o�c�B�� @��P�^���k���L�WF��ݴ�X�{�rC�[�k_0:��+
�)9���(S&����v�D������{���?�<itڐ�i2�{i`@'Ƕ�T>C��j;W�1<����D�2A�v�ƞ���J�)���ln��D�J5�L��J%�C-����θ�I5"���ѯf��x���%U_��Q�{�O\9EՕ)�*�c�LKl܌iX����蔪(סO���q�6���*�I��wsm*���Z�d�ȅ����)�u�J�=�q�;T���H��.���*�s��X��:zyj
̞�O�$�dB
)��K��1�Ag~����-Zqk�x��1D�^��j����.��<��dI������e�\�Nx/M�z��n2�&l��;�������As���Y�������uF�I�}g���]���X�㻤�;�(�LQ>�)*��K6�5@�=��64qo������k��A��d�}Ь��2cf�0W���؇�H�K�������!=EY�ϊ���[f��9�_R�֢O~�/���L��Q�X\���c��5���[i�ޡ䗀�|��QfĂ' �y"̃B5�5�D7�߹�D�ua]H]�)YԶ�~�H��̵�R�A���>�y����G��_4}2�E��������1:�����N���:��̪$�����{}��',0���B��:t|�~f�a����4���s���~�K.UC�­U��
��%�ʫ��s��T�Nl|���62���F��@�ҋf�D�HB��N�� �t�a�^�F��L=5�7a����&Tжf��h�����cQC��
j!���>�B���0߰_$�� � J�	�����s+"Q����^��5bwX).�J�쫵����ʔ��ɟ��:/F�y�-����"�{�~���`dXgЩ��皷�+d�:im�&{R�#��Z���=�Zr/�f�왎���z��.W;d���Jҩtȴ;V�t�����A k�7���!xvOW����~��+9Pr�)���(���m�����B�� QsK�,l����$��\W�ǿ%����4�a�s[5]�����A#c$���9�p�P��XR�f��Ժ�ŦU#֔�n�љ�� �Vgz�������1FON�&=ԕA?RS�'m���Y�e��|v���L�qa�e�+���r\����*�k�����������}M�Rݱz
I�����H��6O�3-(-ˌ
>�7��>�?��5xA�W��F;����L ��j*�V=f1�*g�eh����tO���t9s�����Oo*�h~�+�"��O7b�U�܊�k��CG�<�ʱD//]W# "�îxT^��v��t�����v�X+��I��N�`K; %>��
}��@� ��'a�?e��#�$��]<b[^u>%p�2q0�Z�`�L��5�NWSЎkՂ�~�x���T�hw�ho�\>�C�^��=8�I���W������-�J���'�SͲ�k�f���
��8eS1e�U��4䅛�����Z��4V�.���;���]R]v�]�iH;�o�Ƴ�z���a���V֗Zby�B�"gKJ�������^��E��y��u�TC�N��,�����QvY&�B32��`����3�H��~�K=�I��ݐ-`3kL˕hhu NR��]�O�W>_��g06��b��'���"���2�O���鑷�!��;��
ER�pט1�؜P�X�=��<ǖ���R4{b�?����W��Hh��F�0�qe%A�in��J�)J�J�8@"_�h!r7�X������Q�c[YA�.�D�J���|�d���<��6"��V��p��0I_p�����$ !�E��_��
�_!�v�q�*_�X[Etj!��%���6�ðc{��)x��i�����+Uk�)�=���O3A�ݦ�읐.v�r!�%Z6�as��|�0(���!ц�eѐ�����{�b��]�����t6(Չ�`J��@��&tմ<�w�ڧ��Ńpw�cz|S���G�W�_��|�xtԱ�e�L9)d򊚘���ߴI�j�m��!�22��
��܁S�C�gR{��/pۗ?؛I1;�|���)���;K;�Q.�ҭ���W�˂�PN�/r��(C�n	[�*3�,s&v�1��4�R�����L7��ÿP���������c�
�!Q��(��>}O��&�_^;�h�H7"n5��N<^��bqۂE��otĵ�x�\��b�F��^�}�T�3c�	�Z���R��Ҝ6�����[}��v*�RwƊY"&��Ih��x<�G�"ZdQ��Pʫ|�U�4�%�ڊ��y�q�{K;��K���Y������\�\瀁��(_�	��2���m�y�5&_�3��\\�%v͜��u͂�A�����»^�]��Z�2����a��߫�Ĺ��Mi��'*���΅"�r���� ���n���c��W��E%�W��Nf���������չ�N�c1a�|*�v�7���{� $�Ν�2\ٗ��z����_U��yڦ7����c��өf���gu��PN6M�_�Ě���dSX"�f@`j4��c�O��r*.9��j�<���I	k�M,\�.�뇏�y	�P���T��C�Y?/]%���%�Q�u^|oߊ>d��DOyӄ=Rx�ۀN�TĖ�=���e�j+>9�'
�4e�.h��\3���g�:wF%�@Qr��&T�{,��N�����N��f����gd�Xa�����?��/`���k99n�;Y#�>Pi��X���������D�M��𺐘_�X��;uP�xL��S�,1�!���MM��`�)=�@����h���7�j#�FU��<�A�*�ئ�<�e�eG���Lo߮mG��3�T�bi�~Rq�����Z*���U炢�=*R�a_��p�H�4�/�X-�_F�#��ٟ��3��&�_0���؟��{^���,����6,)ϖ��T��4K�����EH���~#~�sd�6������K਻���V�J"{���ڣG���rthS����T�1�߇qf��~��ulJv5��w�:�w�|+�����9�뾆�����@_�)KR/��9 ⋝42���1N}@\U��dQ-vV��MU��e�{�`�Zs�i��xi�t�3m�F̒N��l_ʉ�����l�t�4�s�Tr�:|��ɳ�IK���Q�,Wp�OZ���bAZ;~���J�@C��Js7�������bƖ�+�]u�<p��F�21�Q�+v�p@��!F��U�X��X�]��d30�Q�2�6#T��Ƌ��Pa�9�@� ���3qaD���:E�O��e:x�n�}�'�A����5;���e�0>���L��,^G��'�,��ƣ��hβ_�ܚ��A=��ȶ�.dub��k��k"l�Pؐ0�i8Tн�T��I�Q�ȧ��T��М�;��N��h`������:�ڔ��F�����v*Dm4�~�z�J��b&*[n?�^�PZ�a��[s�V��#�Ms/��7Y? P9��lo�A��%�q̘�jJ��s���g@F�Y�'����)=��9��"z-NV���;D�����ɔ7�����3��>�d>�OC�4�"��ؔ�D�q�"������i�;b��}��F&�1�0*��0Ǫ�n%�/�������T �LͶ>���E��8����AAE�@.�G�-hŽw>+����4Xh�SF9�8��}w��R�q! ��r9����CHXԦ0�PB�!�WLn�-�M6�rD�!j��L�� _����� v?�"�v0h.�+��-��K�:���G��@G��$�<%[,�e�!,��J��+�R���ʚo�7��s��*��j(�K�!-���2�Ê$�P⾢��mf�)Z�>/�j���M`��j���6h�a���LM;E�l=<Fݯ*�	��BA�q(�d8�C%���L�g�(���Sm��>񗳶���Y�F� $�!;^��|U�D��Eʖ�����5�.�b��(�ACj6E�<��C-�k�?�_`��04@�u��q�������
��dNVt�E��d{�!�[b�ˀ�K��9���wNgڟ/�Cܥ�VDt@���t��*��M�%��@pB����x�l=o׬#k,hc����%y�W�Up�eΣ�5��j�3�,���-wm`����b�"�G1�0��k'F\�9tEA��vQ����׷����M�}�#�����B�v�d���pO�X*�󨼿�0P��О�:�Z��Q-���v��#jz����Co�{-:�CV�6���K��/��UZh��)R�ʅ3�?�4A􄈥(N�
r��}�:�1t.���D���9q.���JvR�셴ؼHn���5����]HH����j��2a��@�eC�.۹���cWg�n�~���g�#��-�$�8�Ε�xhd�u���S�R����L��!r�74���!u����o�/�Z����es�p�|I������,#6�|�g�X�@�W�i����(��h|���L�%������,���օ�vkR��HY�tf����'�1���6~e��!Gu4g�I"ɻ>��e���JFΚ�w��t�����1ro�0ke�U�'���S�?j�)'j�����L�{��aqI'2�� �yYZVL8�&�"��f��>�|n-#a~�ە&N&�>�x���#�_��O��a���=���*�Q�7�1~�	L^2g�x��g���Q��6/�&� �ɀ���`ʇ���`�� �VjA�s0�p����EL��6��}��_�M�{t�Ba������6�@��{�e�"V�m�#T��ĵF��e�D1��E��]�"��6�aL���\��1TEE)ApS��5�<b��.��m#���24��T	�ī(Wڻ��nIsQ{۷�^��p��#���TO���W����VÑ+��1��~:������D�;��*���3�7~�='`��٫���Х�(Ё!�?rvG��K�{��u;�*�O��T��X_ɓF^��hC|F=�`�G�k�c��u�@t��|x�'�@���L!�LJ������	�3Y`T�g<��8랈��q�׷m������}�:J��\51?��g*2��3�Y�9��,��7�j���N�Kg_ff�g����rX"ƽY�\��!���Y#/�[�4�N���zE�Tê�G�t���P�9Ϊ�K�{��r�u~v�G�q�|�Qi��bK�	B�^���q/�ڄP<�50��pꬆ1j�~uMkb�G ��֣G%�d1��)<<�Q�
4�E��C��-�qw��_���SH��A_e��Gy���}�g��e0���e�)��iJ۷ɐX�����
U�;x8��b�0Ԕ�P�a��¦5
�?��sy���A�L�8.�������Y����mPu�Xb�L� �>Ғ��g�r�쏀�[�����7�� �_BF:k~4��D]�a��(��R�v�B�ͻ��4��`�6�^�($�l�hO &Щ��=��O���Pl�t���ql'��14x�& ��i�PR�yr��$)ՠ���+��,RSޡ=�c��m�XZQU9��maly�L��E"�i�F���|����g��7bXD�M$�~_�V�η�<���,.�+��ABד�ԝ����F"�k��k�c�J�(Z0z6�7s��7�?�����D�T7`�f���ؕˤ��2�1��g�F	���yn}L$U��k���j������B�[B�S%m��$*����I�a��oƃhy�c�w�����ǋ�g�v���}gץS����@R�%k!ܘ�>��5��lS'�!�����W�ݛ#�&?�c�-�_�w��y)��M���49SR�� �Rh�V-�q=9À��B�����w��u��GB��oWEb.�A��+[C��/�R� ��ް\4����}d'�dMsB6�����4ۚ�6��)~���.���)3&�e0O��18X�
�s�=�>�?F "�8J"��[���C��V�M!���m5lʙ��u��Ʀ[��Iv\l&���������^Q����4��Ξ��83|H��|I�1���m!\F�DЌ�8l{���桿6H�4D��@���f�¦b"�75��h"F��L�A0�4��}H��j�5�K�d�F�+ԡVC��9�;���
����֖�i|�<bV0��K;S����&��Ų����\�S����������R�0�B�ªJmm�M��H��0#� u���ή���6�;Ҭ$ӟ^f��O�>�Wty=��6�t��S�һf�v��͹^r�q�Y��|�v;��՝ �e�Wǁg^�_Pn!���=X���2i8g�H��l�Bֿ���Sۙ0���#���ir$���ܙd�*T#�\
x��9�e�0�n��A6�g�ľ���yt}���v&�PA�n�-�:c&�A0Om�R�:�>J������x����(G�:�(Jr�5}h�����#$C���3�6�"�E����«��Y�|���Z���B0�rH�U7|�ܬX1�Xȟ���AKA;��a��~F�ڏy��'��*_�M3��.�*�'!�8B�F�k�R NB�׀�S�0�zNX���^m/eR.��LY�%�RA<���k.|MN���Ja��E=�T��J]J�1K��&��#'[�&��@ �����p�ٵf�_]����wx��j�����҆Hho�c�(h��|5,�%����E�`H�h	<�՘�-����F���?�2�'�2���@�N���ŷ�3l�'��S.N�H���Q�/�Bo��g��jc-��%������he��e\T����"G��������ǯ/8�1:qG2k�?\u��w����"�<&R,�dwb�u�!# \��O-;	��(~&D=���ű���!as{Fzƴ�q���n[g�	:sD��H������6)�:կS��W�=����ⷞ"�c�*�����m����s��.Q4~IJA\
2BP1u����)�n~s��3�C�q|gŸ��hlF��F��O� Y*�E;GF��nz)��Ά��d��ݍx��9�04r�#��+
/Z�]��3�b�	�~Q�$��uec����̌D/���/3s/�J��#��9
���	�T|������:ŉ���H8��rڻ����5�}m�&�����{Ɵ�9�w+{��{Z�}^U2�(�&�ًr��x�RJ�6$&���r(����G�.�A$Iu~G?]=�#�D!��sIL�E�M��O�~T�e��;d�ٚ��dVg��7��J9�0�X��.���M"��QA�6C���d;�M�=��[Zi�� DL�^Q��Z$����qvr�ֈ}�aP?�ix$3pi�����a��{���8>�ɂ6��~�,���b�X6?���MC�sL��W,+������8@���6��I�2�Kǀ�`+�B�_�;�r���w���˫&-�,7$����̚<�0��:��7��yX���l��0�o2�4
������Z����6w7�Bqf}���,k �����EdI�^�-&�N�,��!ӵ��# $^�NL��_�pJB�2�ë�FE'�St�u �R=�MDo��"���opY�2=o�K�t}g����J�q��*'�V#x5����e�"�x5��Ka�@l��N���,�Nw�	h��}����9җ��H>u��A����s��`�����q"����*O+�4?X��ل΀�v�+0�g1�$_��(�����I����G+�t�օ.2bڥ��0�l!�Nܤ��3�,qA�mQ�#�bL'�_�|;��Q �uL;�\^�\�Җ�t�x�o��bfY��	BS�t
(�@����&�L���)�&��2	�He&��/k�/��'>^#��?-%޻c{�J����ސ�,����M3�ۨzqXE-���d<}>�4G�&�?���$��#r�%��i� d}nƆ�a	�/-*�i������W����%8"[;4s|��ќg������_�$��Z,�E��8t�N'���%e�Y��aj��g[{��o�<\%�D��I |�$�e�.�C<<�h�3/�x
�VĄ��g���^N�	%���$<�c�&����E���S�G��`W&z��/܉j���gx���i&	D�դf��
cgzpm�^�p�6p�Zq�.XFj�0�c��7�B����H�^�v���tYvqI& �6�zZ���=pSk�;bB�Ƚ�L���ㅦ�3G�~�1N)��!��^.����y:䲵�^�}Πt��D,�#j8j�X�\�W����튡mu�y�(�`Tg06t�`�9�RoL�"|��?%�;�U�l�Y�nVJT����R�,�1h��G��L�^��8$�����+�8�%9����ۭʏ���k!8�D�ƒZ�U 0�<�Q�Ƕ����K<���r�3�'������TW�ٓ���@�e��y� �AR�K��n�����'2��U!EPR�@��޻�I0�ֿ#{/Ű�1�d׼�π��-�|_M��u��Y6������
�pu(<� ����?�R�j����.)zOԮXi��e4��2��k6��i��=p%���<���O�x���8�4� ���;��$Ӵ��;�=�I��o�o
��"�����M�fqO<�`�V&i�+윳�x��!s��/:n,��!�b�����a]�t��n
��Eʟ�b��(	b�� ��V��Q�r�cG!W��6���勀f5��g)�� �AS���״
uСКB&[C����'�s"F2�����#��%e7���xOa����x��aQ�S(\a���O�GG{9wb��\��϶ύ�*��}�+H�h�7 G��(4�&�?0F�䎻��@����O�"�*e�7�6�H����Ԡ5-�/e��Ԕ0�|^D=�P�����;�(`I5�U:+A4m:������ڱ���30�^�F�B�N�+.w��ue��T��\0L���<�ҭ���`� ����V��Z�J�c��dN_���6@��p�Z(}8McF!��)	�؆ŝ��Wv���~ݚ,;!(
��h0�O�(g|��_�z*��-��֊��K�
�t�sK0��X!2����ڙ
4���������SN?�^���W���]֌B��i�/>7�$����3�	�n)E�����}��5�q��J����!*N�����d[�2'q�a�\�I��S�A/^�xz+	�������Ai����(~�����R��2*����t��6<!6�j�N��DVų:�q��[��vR�ut��
���Gh��c�N�^�d�m�ĭ�}�����  �	uA����w57��:Wje챙3� `�ߞ4������Z�0���"g�1"ņ����v2̧g�u:�%�Bb�L�im���q��"��)Ӭ���ْ�x�d���т��߿����w�N�e��i�E��L�.��U��싔��T栮�[[2�� Y!���g�A"!G� 	���ud>�󉣌G�ȇ�7`M�s�G`�{�]^Fg�"�Y�Ԛ%L�A:����5O͕zB[�B���?�),L
��E�v��
�>h���P�z�tX3�|���jwr���,t=��K��I�­~o��U�����F**�e�9�T���Hf���Y(nY�u���˜�҅��{MS�RIZE��w�4S7�u'���-I���n��SҴ�>�F3*l��[=~�z���q�	)�AGnl+yE�tc4��{x��^\ص�)�8���Ǚ�R�^n(&�pi=)����x�pu_�č?P�?	��@�
�"��J��xVҧ��(d�S���u�ǹ��o ��^����=�� n����������;��gK�T�YL�mӧ��˱��܋�~�D6v��n��l���Չ;F�_�Λ̇�~r�7��"�*�/M^�p��! 8m-+j�ts������k�������c��n�χ"cШT��|��A�#�?��|[e!���<F��^����t��|E�"B�%?���#qs�NRk�f�$�1��:�_3�b4��)O;L�I���@�����K���IY/E���Cx���o�w�{�8k�d�~��h��%�H��9OӜ��L�Ƴ�s����2��n��|�VQ�R�J��|����g�3xyUW���m���~ue\�w?M�cں3�̳k{	#����]Hq�{�n���X���h�ƅ;�h~8J^��Ǟ��I�sN�����Զ�OAojk�&sx�I NH�yc5=����Jj%���|o��1	ߌ�*�0,�/�*w1!�EJ�I�0�#7�б�0ܽ���Ǐ���3Ǽr�tˮ��?}/��vFr|>�|6y�N���a0cy}�q� [�d����!�{����21�� �s)^T�3݃oս��_&%�CX��?�B-����^����Y��.-�1��}en��=2�F�X���6�������i`0���9�Z�F�*��\ȣ���bI�R_{�Yi_�Eu��	���@���(��SX��l�T`�[j.�&��I�P��OFf���C�]R�@i�4���Ո���Uwm`%&6��-�vމ��=�SRR�q'2���:Ѧ�V��E���+�S	���h�i���ۜv:/�T���=����ȝ���W �[�V&�����$��ן.���8�ȰU��m�	f$kܫ,�l��&�u���Q��H�R����鰖A��{8�8��&�,��C㡆~[e8��ߍ��ҭ��˻7o y�����#_͹�3�عQ�9�JE��W�\�Pڂ+m��ّŢ��SΣ]o$���ܧ���y�N�X�Be�Q2��jC��?�S�3۬WDi�����Ӹ�	$����L-@<�G�Zh�W?6��7L�H4b�AS�a����r�[Fr[��(!:�m�D�y���p����K�R;�\��d
�}��Ԩ�m� �ƅ}*����n.�*C0�7��8z�5��;. ��vE%Q=��m�0���cYt�Ż0X4T�����Sh!꺂��viQ�����a�c��q|�����soȈ�}۳���t�U��F�o����bBT��U�S�n:��ŘY�!/��T�s�ٌMq�j ��_~K��@jI����g�׸�7�3��^ʍɵPI��q�C��(^0S��J۳kS�z��P�פֿ����j�+O ��p�s�n�<d4��͗�	Ӥ6��踨.�v:"*��Ft��A���m7�hW�3���q撽
gFӕ�x�ތ#��!:�\��O/�#'�r����a�2�O��,�怆�ԗg�o�AV�o����چ�ܑ\Q�Tfߥ#!T�K(�#wn��m�]��i��u k��X������e�����)L�@w��^�6:�a��L93x��=�x%�Ƥ���N�U�������uS�N[C��m;� ś���4e= m���*���+C32�D¨��Hy�l�5o�*�ž�R�@>��9VuD��NxB%�g���!7�M�R��֩K�� {���N֧X;��ք{�E%�b:x����Vvu�(cu���6���~�  ��������A�\ʛ�x(��v-�j�ѱ��#X48���y���.�f��'�/Ԉ&JO�~���U��җ��g5ٗ������%��$��j;�pڪ�� �jn�T�����ɸAL�@s�ktk�谲K	g�S�K��2�P��I/[2��x��xMI{�_FGj�F�=5�.ۡ�>�x�u������J�+�ꁚ���joԋ��q�:�w��Gb@��C���݃�y��H�r[��5��9�!Ӌ�%ҋ��>Fb�<ȡ�ӏ��SRb�ŀ�X�n%h;��N�$z�Y��)��J3K��)�e�/�PAJ� y��X)C����1Kź+�A����v��'k@ꇵ����U�8V��*�����z���p�0T��HA�Zu0To�Nz]�1&Z`�V ���U��Wzmc��x$���R�v��
�x�ΆD�lP��r_���bfN�Ab楐�^Tp#�V:�NV<'gw�~Z|e�O�VY�Dt��{��޻�z�k�޳iL2���2O#�=�/���ߟv�#�#L�����c���d:�Fb;w�Z��W:���3sх.���Nu�I���G�gc�~I`J��w�{2��X�=XBU":i)�Zf���6(�=�y��a�=��uX��%V������e�ŀ9S�����}O;[o��̴��7����q�ae�GM����}Hz��poM��@r0ZO�Q�K���!��Xi�:�L�-��X��5(�[����N9�!1o�y��w�ЊO��VZ�<����o�����:\�^m�A����zSZT�!�5���v��%�^A�\��B����0�7����J��&��2�қ>���8�f)@?���R��n|B�"�E�A�}%,^�D:=MkJqr��=��wv��{�ԃ�˃�~.�@(�\ݏ���3��1�/��/%� �Z���Ϸ��Y���	�7��r���K����A���G���R?SWGS��5�`�;{��A6?�mpӜ�+��̺f��P��@�r��)�J�����;�&{�M�Ѕ �ȧ��7�?�P�K�~>�����(~op���VEp�s�s'Zy����Ė��o��+������{�;�y�b�	�K9��5V�e陪g������>4�M��O���5{����v����#hA����z<*�-�8����f��N	�|��8&_��f��$��[&��n�����[��<����+>�)Q��~����L4E��b��y������m�o��{z�������*�#%/�\�A�P�.= �I���ZZ[+�� :�5�95�,��Z5��۸xR�<��9l�N'���kt�)��NX5����1_%�tH?�E�C�,#u�A��Z櫋t�>}C���u��ڝ���{ks2�߰��%7�4���VW7�����n��F��h^W��h��[H�KY�H�M$�x��Fd��>�qJ�N�:�mp�p��,���� _��>w�R,�6kq���81{�N@�Z3+��g�D��F.�8o|����i�fM6L�\�*���c�HBB�.������"?�s�s���'��qm0o��Ob}D�\KvaB�}쿓�������,�fʑ~��W�pC�DY�R�T�H��3Ø�w��2t��Q��57J�R����2կG��a�mL��?/}xǩxa��έ�]���z)�![��Xn��H��!񕀉 �zd��� �5�C����s��#:9�۩�	�
cy�wGK�b#p"�x�EQ;2ӑ7-e`¶��R�	�Ei�����)�d�zQA
�'e�FOG�C$ρ/F0^#c��������9E��?\���L]vU(!�c���E�4�[B����k�?�R*Q�tbrE_�����`�-y-`���_��a���$�:��'5��Z�A8��j?~�C��<ۤ�s݉�68��l�j�=c��O>�Q�r~Q��
�|ޏ�bW��������r�ʸM������R&����`mpé�+��je1��&#��8�a�R��pwT7Q�,�������+j���\F��9�;��d�d��e2������A@���+����3=��&��yU���[�f��g�����SiF	c�/�X��5�9>w����Z�L)���<�K.eM�ϒ>��BI�"~�,:!kzW�r��=6�*�xJ	����Y�Et �W5��P��j
��+�7{�a���$ fA���2���H���&`� �H(+-�h�'�P�u�������7�t�����W�	,����j���Г�ђ���N��+n|���Ѩ,T+q�`�Z)��Ȟ.��n�n��Bq�Qʚ�\sj�@���L
��n(3ɒ�R��,�b���)�+ſ#D� Ŗ�˰��ڣ�?��-��hM�!�w��{,�#	w��hF���������\7p���D�
�>l��8;�Q��vJF4e{�������FA��:�bGM��4��R MAm��
��[b��6l/P#�U�Q�{ܤ�L��f��[a�I1'"b�����ep&O�V��ɨ��q�u�T��cM3��ɜZnIM��+����:�/vPS�%��Q��B���Q�82�)Ϟ��aI�n��J�=F3sm|3KO�_�x��m���E�=�:��6lfȦ��'�X�z8�AȜ��K�O���c�Q��堗i�B�{��k�X�{�Rj���4$��E�7���i��K���聾����n�����O�?��6�����������v'� (��Fy��pS�>���Z(�F�صc��Y���z����μ�
u~
��j�)��PA��{q��)H؏�c^/C�i�cMnI`����Z��V�1s�Xؐ�ң�ԴBy.e� ����?�j��HU��H���ɥDJx�~�EM�$�U48~�~[Onn�r�c�h�R���S >\������Vٹ]�}C��"�C{sV����2y9X�si�N�*~��x}���0,�V�k|q��KMl���]����#�@�[��zñzL�N���;�ה�O� _I%Gӫ�:�����S���D�$A�=�L V�����]��l ���K����d�k���b�H`���9��/�(��C�l������R6b�BC)~~��Uk���Ʌ,ld��~U.�A��fń?�j�jPDI��y�6[T������I\�;F}��=�L��3������3����|��C��jK��:m�3��<��<��Z!���Ɏ�m���z�}0�8+�8���nv��C��|*&,�0�,;G�x����u����"�)=$�\s���A	�
�Q����2pu^\r���
�*����+zW� �C����9M��b��_dQX}L���E%f%]�˛��ס,�3[�b�s�L���*��g����� �)��{��Z�Դ���2��=�-d�叜]ю.G8�n����S]4�rP��F]���Tr����ɋ~��a�Y����v�	���R������$�@9�Tbtq�^�"��I�Ay�
rÍ!��z���Q�w)7(�V��t�O�$RP�4��.��5엌7� ��s�
�:s��p��&>x|)	�_�~�<s9Kc�u[#LRƋRJ+��Y�7��D�U���,	��G�\x�f��.���ޜ������>)�J>g\��<��l�����Q��2�B3�"����h��
$(��s/��8R�9S��'���z�OyM�Gb���e	�E�U��D8n!E����֢�\k�V�"�D�?U�'RPF�����b����S�ٍ��$#���Z�L��ȃ�^�j�є�ؔ��θv"�0�0�V����(#�� ҰJ�m����ち���Le�ɺ�(,?�����1�/��̖�0s	n�@!d�ᶫze�4��}��S��I܊����(�-ކ � 'o�,V3p$�������ݴ�b0+�[��" ���Z4�N���;�.�˨�|!W�C>��-ӿg6�J��j��Ɏ.������������a�slp`rf�>5)��3�P�:2�J����F4�״��I�JF��S��P.�Q3ћ�����1
�܉p,+4+�`���e��CE�,~�kj�S1�G�������R����f-nB�;�������g}Ő-?C�i��\u�����د�FX�!�V��Mp��#���9�4�+��z�o�F�	?ԙ��6�2M�_u��[�!���ٶ@u<˦8��-��r���O6i_,�%\Hh�@���b����}��7�Þ�q�V�j��2!���f���ˀO��:e��=��0���J�[�F��nC�*h�c $��H�{�B+2�Z�F�{F3�!��y �0/w|�7�Ղ�.�z.!)V�?�qcY����{�!H�&���M�B[덤 �{�+�/|��V�-��-�-s��g�1 "Q���hAL��'&<@uͅ���CpS��M]�(#�ϯ՚�/Ac����d�>`���:��(/�#ʰO�����L��v�xs3��T��\�W��JM]�R䨐2��0�٪�GZ��r��X+7���%�XQ$�@���,X��e`�Ps�����Q��Mw�Gy��Z�we�"$�&⚶�p�{�a��,
v�ͪٙG��kC�ԏ������Y�\E������=���[��pE�Q����~�)-��qs�n��/&���⻩Р���Qܧ�mty	�=�YQ2`��5�v�vJ�����F�9�A�ʽ�A���!E����a����!�R�Pg�� M+#�S�ח���~j�T��ͮ7h�~�?�ܰ�vO��a�[>s�/~y�K�#E�&��Wx}�o}|*�v�s����9d�I�1{��y�9 �ʵ�r���`l����,�d���`S�����L;ȇ�$R2�䬃�
/�7�;��!X��/eQ �4�`�SE���c��	���l�}ʪ\�ti�W������,�V��؏�%���a�F��7�at�}Qc��o���{ ���߭z{
�A�Q����������)�y=qό����:sru��H�4��}rҨ��٣��b�u����x�n!tA���"~�3(�l�^�`/����\�7��|��#�n[�S��Й��l�$8�4>�`�d��B쥄�!�ߜ�_ȷ\�aB�1� "X�|&�V�%�~])�b��>�9l~(c<�kZ�Օ���M/M�;eMTU0����F�@�Ix�.�ؙ�M�>��[#&��j뀚�*]�y��u��Z�iœ��u`������$(�͡,�l�ԋ�T�J�gž���Rq*O�	|3��q�hTH���u��=�����4�nx
�CJ �����Cf�������n�s���I�z���O�_��M��|�O�c��`��������/q�٢�R�'w����AH����WW��(���a
�z?u�� Q쐉����֫2ׯ���b�e~C�N!zT؀���[ک��PR�:ڿ��;��R"�s�A�N��o�ɗ����ݏ�Α�lBd��;K$�'������p�K�c�T�CK��,������'��1�d�'i?(��P����q�ӒgG8Bg�/l'z��^K���V�\A �RD�E��gȄ������m~�Ȓ]ۍ�7���r��~���)Ji�A���$j)E����Ҷ��YC�4/����j��aY{D���H\���0L���ݲ�F ݟ+<g�7�ڎ@�&v[g?��g�P�mH�nsKy����B�R-?7t��OaKc7 �vkJ�I$-��\Jz��+��Q���PV�V��~~xe (\~��dc}Ue��̯�U+�6���O14֕��4:�����L���Ćn���1�,��\�✈mݿ.��"ݶW��T;�1���;�sY���nϛ�2N�Ew5�
���� �g������K��F �#�N�[ʋ�gr�Q���DEȕ������p�JR�Q��V���Hu��T������j��5h���S����v��Z�E�s��*>�q<Ȩ ��5�wT��d�X(	4{��ha���
0��SX�jA	؛�l:�=@mt����`2O.r4��F����Ev=�j�yt��*,�?̒�UP��]�����>c���Nϊj;	S�5�4q~�y�0&_[o9�):��Z�[X�u!=����R&�jY��(`���1�gu���g4�-P���R���ސ�BM�1���thL������Ȇ���?�-UOL(����	s[ߎ�'��_xb����sq�ܶ�� �^J�6��Ce�
��S�Q.(k|�ΰȏ��?�e�	vٱ�{�	��_(��30��!Q��1�M%�<K]^��U������|�ꥆYNO���	��m��+�]��߂�ڹV㛎�fz��З�T?�*�ĒN��{jyЋ�no���'g4)@�9?"���3�2�Lx���f�YӺ�
`Wչ��gn�J>@B��|�m/�l�R����<T�ˣ�cx#b�
���ۭ*m`�K,��.�ں�v�U��|�Q�9���� R�.S�v��4�b�@��aL6Sd�W���F(S!��P���-���9|�M!xFK:�Ѵ�/�����}�/��S@S�&fj4>����يz�|�>���xB�dc�1h���z�l/�_}����f�p��.�J�R�s�_�ț2��:�6��6G��s�~���6��Q��� �::�ē�q�QT��������:p�d�S*b=ަ�rN'�T)���Ƞ�B���k�%ǆ�s��l��(�d1��z�x�b5�DMv��ƐeZ��̶�֓�8��JH�8�fQb�zo�*��&ӂ$B���1�$��C�>3@ Rf(�����8��<�g�3�*Fֵ�ͭ���z���Y˩��ڠ��C�#��?��� �Y�Ǝ�*���� I+*hܝ:��p��;ќcl^	P ��B�Ԇ/����`����L_t�@���m�i]�)6����=���W0|XBG����m���wvo�i)�����#M��KoK� ����O�g!	��솄�)�����.���[��3�f��i��qƹ�����9����n�����R(fk $���Ȏ���'�Qm~��C0*Ee��� U����Up��w���1��l��lQ@�ܠ��\ͦS%z!��=��o<��^�?K���<u�V��I{�)N1���ʑ��5E��Yl/u>Hb��o%(U.��C��r�a73������|��������6��T8�C[#�!�T-����P���,�r{)88�K�{��낂^�7(�&Rr���\���/��bg�7�W���I�\<�$&̀��$�0Ǎ$O޺E���Y� ����ڣI�R+`^a�	d��$nG�m �Gc���-J201�K�䃩�g�v��&�����A*y��V-�@�X�^�V:���АF����O�:BoCm2�+h#jfc�
n�o2r~���S0pJ��g뎒�����N]ކ�)�-���A�~슓����z#�ڷ��CJ��u�q����t��ׅV�&��8���	h_s�n�Iu��*��H�`�g����t�36�h���s�]�Z}��ؕ��Ԥ�o�˷Ӿ��v
\Z��S|�_kB̎}I�W;�VOb��7���(X_����������"�4	�D �Rq͞�$��>x�r
��dG���x`zUV8���n�/�es�r�o�0j��@��ܷ��]8��)@G/�/Zzm���-��pkoG�ZZ����0l�Q�9�@�I箵����#�m5]Rw�0�i3i��uz*3�L7\.gr�n�A�y�"����������(�4X�'�UC$՞��W����Cix�^��>�jg������=�M�@�F�eG_�j�#~j�T����Jrj��v�?�å����n�b�l�.�SZ��-����s�� r;⢮]���?Ss������.[�_D�qD6���Fu����H�H?�ݕ'(��ˊM�`�$�H���L�w�JC�F�M ΅��6�	i���=}OF�#����eҪhI��,��(Cd]H�i�5C�]V2�r�����]W�� �㚾������jS[O[j�,�Vn���jܵ��=�n���H9���7F�9��6���-�GFEK��D�l����NzN����b�U���X��Ǭ!��2k�E~�z�K��񧐄B�MUz(t&j�Z]B�}㔊�2��������!w�ۼi�A�;e�uR�Ỳ�ds�U����[��T݀�J���g�Ȥ��n��|�~(�,.�OG2��UG���a�6<w���P���Zvoh�T��>�2��o�P�P���qe�jeK
��d��{I�Z4S��6]˺#>&�	�� ���$$��C�[�z9��[�n9�
M� ��
WX(N�{l�x�[5�R<R���$(L5}ٍ^� �D�G��Mp	�7/pƧ���9���i/ƭ�Ѭ�Ho3B�����
ʝ6
�)�I��&��=L�0.��e��|����H��+k9_E��p��?�f��札o �ah3��.ƭ� xZ+ BT�yք���.����]��
�����Z��(�d����4��Kb���OБl=��������L�E��h>���VPvF��,҇����4�cתL
�y��	�xc ��\��lx�}�`�A�>����V��C4n��]CQ�:�or$�|Y��k5��j)��*���R���2�`�i�m�a_I<�*x(���IC����ː�Ż��y;e䚣r���#,��*Q�`;��-$��_RXR���g�4�<���c�w%�����_�sԓg <F�6������~ъH���d0W�P-���,��',)hx�,��%u�[}?�б��c��o�T�3��"96n���|�4Ü��(���Ik�l&Pt��N8�=�CĤ@���c�b0��Zġ��uL��K�
���0w����i���������:��:���,�M�W���q*)�v5>�[p[P��9������V��m�����`n2'r�봡�bޫm�1��)���Q�5X�$�8�Ū�?�xE�'�6�����iI��s�s�!�T׊��©��Lʹaۻ��J�%��0H�윤f�����J�ic]��������E�1�7��V-����;c9���XOR8n�ge�XǟeL�������
O]��^Y��%�����H��>��P%�ȋ2�$)#F��e��	x����Lx��$o�5r��[S��4\,�/�c
H�����q����یQ`���Į_����XXݭ��j�سW�T[z��|&$X��{���>�S�����d@)= �ڨQ���V����KW-ޛ�e��Y���ޞC<S/�ż�zw���/�&��-�e���̌'�i�U�	�g tP�����0��M�g�CE`��D½&=]�eb�a}���T�G>h����o2J�����]�:-� K�_�F�\�6��ϱ��u�`L�����QӛM5�'�_7� �$I�f)�������OթM���r.�I�X�P�̓$�煣��Mci޸�M`)�!c�ǎ���Ch�pj�")�x�E���χwދ�g�+;��R^[�L�苙i�Q��1r�{l�G;gB���9?d��*(*�H��/"�p�����Qj��@����;�<�f�!�(R K���4��AS���0��� '}�G�a�X�K�0�*`3���
Hh:m��]��Bʞ_�1����ƒ4�����M{^'�k/|eR�9�n�"�낒�^�Lfn�Qʳ��A�#v��|�ԫ��2SA���${%I/f�Ã:D��

�R�4/�#f�Q�c��&��]��,4r�g�밹{�lȴr-�A���r+��\Ό�a��=�
�~�o��)���đ��� �>�N�Y�����z������p�q�^��苅]��?��Cn ��[���V �g��6�lR£^:�.��I��Zէi���ZȬ�1�f��d3"�Ki-��_nKoxD�M�(c1����J�Zl��6qA���OI��y[آ,�w�b����A��H��	�E�I��E��$��D+�Ѩ�#�vc�mO?S��[	��
���X��@펥h����p�y���+dǶ�x���$��e���e7��hϑ
� �*����^%��j��Oa����R0B'� ��e�)p�8����D��ԙ�/F'�߽�bW=��ʘP6Ptx��~�Nã�k�sYl1m->�����BjIWAk"󞂃��`��an0�x˿УIG�y��j�8�6�e�h7�/�����=(��ˢ��$�2M2��3�=��YOF��d�G]�?���t��nB(�#��)�����Ϣ�N����5|�	Vͽ�xƗ��0��T����2�k�ԭm����/mx���F��Y�f���v��:�W����19_OhUXn@Jh�Hk	J�A�P@�T���[=��K�rLs�b
��%�ݺ!�I2�Wf�E.��.@��F7r�P�EӵlL��|�c�R�q2V����5RY24 ��.'�,W����ė�R���ew��Al��qz�~ڧ�I,=ONA'��{]z�,�?�0bDLU���+PF��Ǳ[*U,O!�I@tn�Vai����bֽ�L����(#`�X��*Ѿ�YX3����b[�ˆ�`Y��Uu����u%<!sC>sR�M�uh�N2�BI֚q�ذ
�a��%^��NSV ��L�@���SϏ\�&�zZ�71	�^ղ��Ml?㻦�\��������q�;7��(6a7CZQ6u���W�z��a`~M+@����督�I�6q����z����۝	g���?��� �<� "K-��1�%b�b7�X�nb�E��h�y@��*6,��R[�V}"Q��I+�$�����r��~�KF��g��%vD9�������^D�2˗�Kx���~ǫR�(&}�78������~���p�`�w�5��<�>�h��(4���b
���; 1���i�lp2�ɠ�	��)����r�:�wv8MF���_��޴P�Q>�w'3��l�&�D�V6��,P�~�!��Z:S�5U$ǂ��:8�ݗ2`�!��]'�,@086��
 �X#r������c��g�Wכg���4��N��z�J�u�1�\"�[�e�/��Ǻ+{
Q�<Hm�:�S_���#V�t�%�f*(�O��ej�B�L;�c�/j�PGI�y�T4�k;�7rh�+Z_�7^��A�/JlnSe�ElK�%f�l�B��}��o'p�F�as�=�Xr>w�m&��	�� �UΟ����G�j�S�+��/��}k/g.����偗�m%�� �z�yC�5��e���R��xz�B�����Q��μ�?�.mS��#>"�����/U4�E��v��Ϻ�� ��o'��p�,4� YJ)��tW#��)���e�NV���K�S��J�GGy:�.m�m�F���FeSu@jʢ�0���7{J�_#~�e�B.K�w�V�-�`pU�D���>U$U|&Ǘ|2"��&L�v�aсjZ�1Ek/Y�q��4���_��X�@ӊ{㕟[7�&�h��|��� �ǱG�m]o���|�.�޾����n��Q��E5���:�!�;�b,]�Y���L��9�GƝ|4����|�#����zjȀZ��/��D�#⏏�N^��D��Kʧ
U����{~M���3t��H�#im���c�@w'9bx�&�ba�'tȴw֛F)#����"�7���f����`(�/�����뗷qݜh+�����V�p�a�c�'iZ<UF��ս��*t��	_:+[WW1�K��bz�?t��a�JY�V�SJ:�k�%G�S�9��b=QFM^IS1�ma=x�V*�����>[R��6���*�����AwY����jO<@��	���Rgo��MW}��~�A�n:�{�M+A�qW���
���;�:/�,��_��Jo�X{�<Y��B�]���#�^ګ�P������*����+�5�W���	G.��U���k'�*&G�vzh��qI�����랛I�F>[A����#�_K:���rt��I�% �ڼ��W��[Gx9!��?������{'tم�2BS("&BDqq�DXx0s"�U�'F�ӆ�x�^�1��Z�5"��y�/
��e�)��ؘۯƾU�nZ� ����+;K�*��� 9�y�y5ݲl#�{f���V�q�N�C� ��nM�?�l�vM�/�Xz���V��J�I�nWҏ��k���S%)࿧�$�u����vZ'�\��R���YU�XE9kHٿ�9W�c\�����>[C���N3 �X+ˊ���瓬@�F]t��w�6�C�/Sp~�z\�)5���b�+,�0%L(�І������G��%u����O���R�����XG3�,����g�{9\�>?���AM��u"��k�dk��q��NSז�����]��1�����/�����~6��|O!w��~Xm;��P�c2WV���:����X�k"<��5�W,���B�~K�H��BՉPF����eS����v�PQ�$q6�!��5�����ɗ� >R9ՃS������P�32X`�7�"�e��;���'�{`�<)�MC��t��Pgz�}u~C􈂌���#^���9 $YA��d�: ��Uo ��I=%���׷�����I6b;�-���ަkܾ:��Hn�&�^ڕ���6�x�Lceo��{jDPH���'��/��D-j�V�g�r"�������b�#eތl}d���,爉�u\Y�:g̀lHK�,���?_J)oE'f4��0��>[_B�W�1��"��A��kIH��dm�Mu�4�!��\ߌ���y�I�Ϗk�����@>�1�\�V�2�ȫ�<~_�o<vp�$�t>�׹�D�̆�M����6�>��L��qxm�[��K����Q=Еu�3GF:��D���ǡ��%�-s�Y"�TuU����ͮ&���1>�ts�� ��h�&30��nx�2�Y���M�,�cO�z_jHY�G`�r�A�ubH��N�G�)��T^��V]�(�ī� ��(���)Tw��k�13�w�������"G��<��<{-��N�+�7����*�Cyr��_������nQn��\.���-�{z��� k����;z���s�&;O��]yG8n�i`~f7F�"��ՙo��.�r@��O<�DC~����8���{���yt?��!�$i���rA�-�:2�pPpd�"�?��}r��G����&`8�[(QLm_��,aw�R�E�|`)��m��^b	oڅ�o`DfXu6�����G�+fKzD*ThFN� ��y,��m��j�@�#0�wWY,��&,!�b�Ye�6��B��y��Z����1~·�k{���;��dNT��i;�$-��T qc�؀.W|0�ڳ���+�h!�C��R�n�g�a���/��v�&��?`A�u�$%1�8�zٵ�Lv�]Eqr�c�(p� z%Y�Fmd�%����O�R
��6�t�}�H���H
g�1Ѽ~��ꌯr,��3�|��+�O�7Q�M �__	��I���o�ԇ#u+���j3��>I�J�ő��8�9z~��?����A+N�ŏsEŃ$t%�Cm��9��1�T�m���'7���h.�G��V([�_8�N��~�Q(�)�1�.�T�RAT1egv8v6Ǔ�~ ,���r7<x+��v2�n�M��1�Q�]g!Ɓ�����b�X�Rkh=�5n���g�=�t�Q�%c��{����q�9� ������hK-��Vq�p��!�p4��?iM���e4��8^���#�žX�N|�v`?�t=�Z�"�@��E�}��O(�ݪ�}=O�)7�M"�K�;��d�y�)G���}��#������V���F�� �m[��
���eC��7-�6�۲RIv�|Կ�e�e����p�� ��m �W���bl|�lւ�0��Uu�0�-d�!L>�tW;`�q���m���j�\L�<H�(2�n�t��8#���<]���a��| ���Ņb��Y楑���hO��C1��{h�B�A�b�>�R����+3@i��ڜy-�k�s��v9����Uy��\�{M����X�O��ʮeW_���,�!!���~�_�
���L���V�8�ǀ�h.ǂ�ܖo 	Ȓ��(.��4��MD*�GR8��'0ی-��"����uÂ(٘�!I��7�
�h�"��&�c�GE~���)O�@�4�9�j���{|pH/lN0Cs�fq��0��\	c�G%��>6���Sg��{aN���U
��9����T�2-n�y��ˁq�z	��L�w�K�1�������B���\o���2��,	-���-��??��l���+,$w�x٫-?U^U�1�H�����] >����eU��3�0Qa��K�WQ���*yN�Q�Ǔ*r�l�<�Ӡ�E�.t1v 8�%��#� V��x�.L�9"t\ߏm���]W���_L6��Mm4nJ�(����+<�
'r�$��p 3���*^M�~E#1���2&�V�a0����g<��tVr.HSoh@k���n�M��!ʌ�M��V�a�4#q��d%R1��Ά�jo������0:����#@�P甮N�b� \J_bO�Y�
c(�պ'��9�*N��v��N�B�"Gu,��x��]=��"\d�Aּ`-���/�B"@½�*P�=�;ˠ�H
���XPq;�Z`����0�י�j��4��,��w����2g9Vd]��j_�b�kguC��z�U��#y�Rn9����-��_���r��! ���G�5{��S�@���˪�s>)�2������G��?� 4�/X1�dCz�5G��PL�Y�Ǜh崵N��^�H q�ؒ�*�l<�����;���O�i!�П��Zw� �,A���h|9���F���펰�0gF]ݝ7F����,���Z�`� ����/1�.�v��k~0T�e�g?K����[����]k$E�?w�?T��Ѹ@��I\���4i�ct�?V��3�\��� nF��ǻ�����f��A�8��T	����&um4�Й.f(��S���i��%��/���H�O�ߨ~�L*��eOT^�|�j��0y��!Ýv�_�IA.a��u��3cgZl������ͳ�ε	�qT�f����M�%��f�Σ#��q� 1��3�`�y���R�/�^�Z�J0Gu����tYw�/�r���U�/�뗜��@@��K��p��vu�C3�ߋܹ��\Z��љm�#E�cZ�0�آS_��	�XV�~����U�x�GsS,*�Xj4�h��	D�g�̊ԙ�����}[�������a[�֨�_n�E"ڐ{�m;U*9���TQ
���Q ��3�%��
��5�y-�o3��0�F�I��̓��4tP��r+�67B�_��dq�tG���0��T��c��!�d�0fD����݌�w8�v����9�c߸�p�I��8��OX��w"��`j�䳘g8�#O�QI��J��\Ww��PKZ�c��8�� �J��L�W�Y�Aۗf���1O��=q����N��H�o8�oP��WP0�Ӂ���+�R5d���������?�f��|s�0F��k�S`�$��]y��3t��
"��U��#��t]XѪ1�nf��A٣�=��*Qaők��i�o40a�v�%f��Tf!^��Է�5��P��A �o�|/����I������^���re�F3���"�4M @��ؿIfc��K���,q���6��OK���	�V��d�M�u�u�N`��d=s�{l��W~�:?�AE�j2��j����q9#���B-�EϤ�6��aȰ�{�.?�l��P�C80Ee�v̤8�eYR�~�!xiי�||�P����V�=��ĥOS%��Ѓl�VV̩�	��?CK��D��t��+=��F~�ڋ����1�����5D{��.�̃8�`��eB��j�,=��N���ow�͊36yt����K	r�|�yQ�ʆ�6�̀�3��S��?ns��>;_�����E$˚���Һ}�������K.�!�;��z-��<��w���;��a���1���Х,x��$�Q�=G05���"I�5���k�\sG["|�%�ឣj���w;�j�CK��x\���ː4�tV���ҹ'�|{@u5
T�d�<I���I��劀�D����ad��}��f� �i2��z�"c��W��W<�%k�����=�QE��2e����>^�����n�9�@�!��?��db��"$�e	RKpF��0~���}|c�R��ێq� �.���D��go�(=�@m�ʎ��:v�� >��O$׿�e��܇˥ʎ-�֦$�2���h���5&�c���HA���y(`��Ԥ�C��0w��˜>�w�7N��>c#j��k����Y�As�z���ջ�a1�T�^�#	��
ݸ��1�!D�uoaK�V����v�1�]w4c%��G�FA���W0+G�	�����.[���퀋��A?�� ���:
m��um1AĲx�.�W���ۄ�!f#�f��dG�3Q�`��B�ذ͈�a��T&b��;?����qNAf���v�FA�KPC���/遏�Måb���x��摡8�8��ƻ���)�E�Y��̚��,���3��'�$_����D�1�m�$��*���L��/��Q���^�3
�챑�X�,�D,]�!�xt�0Pm�jo��ah�	?��"ۍ��pp��5P`���1�[z����;W�j��������V ܢs����V[l��xO�,��J�Q�z��]��5�ó����"�[��E�'��?� ��������jS}�?��P""�b�D��!w)/uJIS����巒NM�wNڵ�&���f���I���YDC^����v��u��}G��?~�v��	rx�ϥe���4���_��b���W:�\�������&���N� �� Ә�|� K�(�Y� �صŬ�;�,�����<�R2ŝ��>I5��$���mXQԑ'1
q��t�՝�i*ң��;�]�n����`�L���r�',���?���x�S}���C�	,2W���S2x��h
�Z�ҿ{��>�9�yn�T�."_Y�j�aТ��4�7S�}�m�nM����Wm�5b@��#Y�H�Ͽ��l���Dq0%C/�� �TjQI��t����Ӟ�"�?n�$�-؈u�R��~ �E6Q�U����9
�GO�~k66�a���/��qU]�>��sg�1}�k�K��� ����w��[AͰ���� Q�����?�k�N���t�]��x�ɅJ��o��`<������8�&JI�a1�,p��gz,���X�盉��kCh"c��=���jM���Y��c8g�c+�g���y�L�_�&��6�����t���q��b_����\8��=�������0r�:�o��s�L�y"{
mg7|e��7c����͵w<w�ނ`'�Ң
^���l�-�\Ņ�c��ù�l���ވl���F��3���3P��.��ӽn�:�C�����_y�ӻoVYx[��s.׺NwQ�����a�X�< �6E�k*���
�
m��� xKRYg�5T�DTK��#�7oW�|�3���.m��ޑ<#�^�8��u��W!��"��
�ea��#|�g��E_���������Dó�&Ih�!��p.�J3��������ö�/L���_@���O�kvu����2T���G?U�/,#A��ܠ�P���ըM_w]�M?�3�٭�Fb�U
:2T ��u
��#�*�b��86DY|������u�Ch�<"��PJ��VA�2�˶2�ۇր�o�4cE���?�D@��Z��}��_8�z�y_��U/�@�{�\SWr�$��04)������]�b�&�{A���Xɹ����Z�4���C�y�l� ��A�����
Yb)_������s0�@��>U:G^DM�!J�T�����O���;�e���R���|��R��,}jt�ᗕ�MUt�D9,���̥�����vZl������H�:��A����Q��T���id]�r���i�s���:�j�+��5p��*W{�x����tȟ[��u=���QA��t$����斟�N�_G4��A�9�\��:�y�[ZoA/�-K����NQ�����A
�֬��ƴ�J�&~D<�wg�f�b5�RlG�S�J�g���7�{F������u<t�O>f��)����U�D��~Q���.������F��B��&�h��>�j�Kz�:��S�-ʕ��r|6����11�w�k�E��i��:�a �Ӎ*�X~���%�vf�0L3�ZK�1Zp��!϶��b���-#���\�wS4ɚ�3a��D3!�m�:��f�����]l��/����6������zoAA��3 <��벸����~����6TE�
ί-{^w""�_�����n�{�Gy���zd�M�,�[�cT��d ���Z�����P�� 1��Np�Ț�3��p�pOU����-�"��;�}�`�/\����ݷ=.u�;u��ח?Yy�k���`�ZֿI7�taU��P�Y<`�U�A��}���˶�}�4?����:^l��z��w� P�O`4�2�&y�K�sK|l���� sJ�hb�E���{(�0T%�`ji�I@���z��BZ��ɻ��Dj�*~�څF6�D;��� �iٴ���s��Ϳ�7�!5z�j��c^�������X,r|n��#��U�a�!�a���</Y*��	���S�~�S� r�{��>�d�}���p�B��'�\��JPT���!6>p_'<WOX�MVt�0�[Kd1����$dN���;>�dAX�0Q��@�e��� � ['
1�y?N����N+c8�T>\�(<���÷=�6�ᐮ��Ow�L��}���$��?���O!"�~f?�Lk9%����73�8��QO�^k�ۘi�-ȟ|��]�u����ĉ{$�K����rjm!�2Ռn��E	�W��{G#nx�y땳ї�,�~�MOX�q���f5�� �kO_m���d��;�����6�8�`wg�>�J�'g��Y:sp�-&	���w�\�1.��Z���Ў���~�@(N��`�A��P��9婇�!��q=k����W�S���pl#dC%���@�H>�R:	A��&v�����'��V#}-?�}���1�!�v��~��sg<�Fx"GoߛaF��5��-���k�S�m��*���
�v�F<��ũ���|Ǩ����(��"����~��
5��%����&e>��u��x���[}5�19���m�Mu+�g�e;^%D��@Q��u~���zU��	韆�7�N�.
�h[�@mj�J�{�P��׽�{�خ{r>�O��|�i�-�]�%|���a��$�de�/�����x;��5܏T���+[_[V��Z�~��9�*	f��8#�Ϡ
��%��(���*�3�����F�V&���~t�*=A!BQ4kT�#�]�L '��`	/�s�������A��
�Ʈ��HN~��� ~�+�Pz�a�Ӯ79���e��C���&s+�>ID��{�%A3�B��8e%3T%�*�ӂ�:�����]�9��t�x�n�y�ݗ���#��R��[rb�ޘ�O��(gv;n��K��r�?Ѵsx����$>�����Gv����3�/��a3��⏹�:K�1�:���Xf��ʟ17�t���Y�{ǆa�j�@����M�S/w.��V(*��b�n�#C���������QÆ$��u%Z�[���t��}�<*UC�}��
/|��b!���g���j��+c(�WC��a�>�a� w&{]l���NF��-��laM�7>��`8{EV�ٽ-#�.�Y��3�JJD��*�%w ��轾hTG��6e��M���C��:r�B����\�a�_k�C��_�\b��6{ѽd�8�>''�ȮC*I�����G���_���z���v2*�+���[��O�Ho���kp�E�/
�Bu�Y�n����K̗�`;��T-�9!Jr�ǡ�/R�T۞��D/S�`�c;�ъ9s �D�xh��xs�Sui ;���9���D��r��� 1�h��j��;����4�{�r�5>�Y�ډ��`3&wL�]����I&�x��#�����18K�R�x�������v�����������):�p ��p(G��4.�����>"g��neO1��C�k�E���-�Z�A߆����&nZ'���vMmp�G��@�F3%E3(+br�
LX��i\�h-�6�s�Uc⊇'�����Y�pǴD$�\<d��^��+���r��ˌ��#�܌c�n�'��M� /V%i�R��0"\��_���>WF{��S?���EC�Ic�'v����%'{�*����D�H�yЫ��S{#H4.]ⲩbqo4o����w	ϓ�,�Q K��:h}~�1N��4�� c�A�?GW��H ��2psz�Fu=�n��Z���">%7��c�$�<��2`��-�dO��9_fh�s�QI/p��� ���6�A=�����NENݖ�_�M�)�Hq�C�
}X�F����KN�J�V�H�~S�潸�5dw�������n���b����q<�ỳ�� C�ɾO��M�Tq;�������9v���%~3.��>�����,wG�� "�
��k^ճS!I�W�?�e�ע���Vm�B;H<��_��ݵ������k��`����Pv�����w'j����H�J�h��|�q	�n�Ě
�t��(�nM쾪��_��_
fBt2�e��o��,S����7��Vw�!�`��Emt�N�����kb^Zq�S��Q�{�ϥ��������}EBe�F��"#U됉�r6�U�4���ɫ��I����3b��I�H|�N9�
=jQ�R����V�3B6f��KLI
F��Ř�w��o>k�ۻOa���徟\�6�v��`��k͗eʣ�-���T=z&�L��D���� +E"�#b���aH�y����o{	>����i=Lĵ�+Wl��3����&���5�U��+P*�!���ו"�I�r��Kb�(^��f�7䛷�W+�%���>t�Y�J�}�^����`a
� �3��#İ�ޙY����7�P�ƨ�}p���mQ�����Z��t"��7o�7/�����\*Mg>6�K[kB��}׈��WMY�p�7g=f���Ӟ�5�*­�w1"�卥p�<���\�b0.�iR�V:|
���b7b=AÒ�o�?���Z}�8�����z�Ԟ�aSX��λz�p�ݜqP�[�yWR�#pN��EZf�~�T���c�����uq-�a���f���'iw4��"*�+�Cbюn�O�
�&
��}�G�-h%)ͪ�vj؎�IM+Z}mw��0�E��@�P�h��	���E���0P�F����(���~��2�⒕ټ��/%_t�#�%�;` <��kMQ��hN�wV�?��l��4%5�^-��C�~uwcD�.�l��?%"aP��/��Q*D��:x��!�OB�s�2_��j�H��a�d�No�n��-'��=�~椖�0��RTn[�l�
9��������ڹ��x�{*���B�2`�]��i%;� �=�u���O���gX��)z�{���x���՟�r�n��}wx�k&�,d)q�	k����.J<O�u�g�Ia�0��h���8�=�ʈr1й|�A�V�lG,���FR�"@��X��l�M��I�G�)^���r����*���w�ʢ�v^F�6�Г�X�Kzeڊx�)-+�r�Rx���d4�Ǭ�E��=Gּ�B���#:����fnC=���W$����( ���0")rp���7'.��RXOƃ��?��'8λy���ș?楿48ݍ�6M!n{�nc�	pY	[�/�*�.�B�N�s�A_D��}t0��ݰ�K�_@�S"�s��/��&Me�ٴ��Zpw�C�CE����A��<�����XN���n+_
QVW�K0���Hv�=�I{h..�| ��}����;�T���=j=�Xǭ��f�b~���v�:7����iS�;�� ���rc'K���_󘉡?�}H�t�|Z��ǳ�M,ЂX���c�!�|Giƴ��3���Q�T�{R��W�d��P��Qbw9��I�P*u��!�W{��|Q#����:��'�����M�'Q%hv�dD��2=��yT���l�I�08�|���<[߸�N}��#����y�N���_K��Q82`t���?㓫��;�1xw5
LhưH�8bh2��&�G���7j������i�L��,�Az-!�
?��++����S��V��L+@�j�C���H��v�l@VҔ;�č�ԡۈ)�a��.�]&I��єF6� ���/ �C�����՟Em1����N�,�b�<��dX�,d�?«ŠwY�P����A!7ӕ�Z@Wܡߑ5ը�Z=���,֫7g�SX?A:H��_P�u�7���El����s��X�O	���l4o@I'	��5,�嘞Të�tI	(��� ���lZI$��;���̪v���)py^��#�6񦧹� �>��`�O}�H�
��_?*�9̥�X�xA�_=��$�#>͵�'��t����yZ���_�q�.ڴ���EHo[I��]Ǿr�}�[R�ף.�a������/�Y:oP�Q��q�})��q�[�ŝ�e��^um��D%I��Qx�#�¸�b��G�t1��L�'�4�9%]c÷ڼyI��x���7�M�
������`�A,՟��{M�$(h�>�*"�]}����wV|��-�O��W��ZO*}'��f�<���}/Έ��Ʌ���u#E=�%��Gc�Td U\��ðf�$ �v���l�1z0{�p���5�jtO�E�-�����^�*ӵ���k��C�hiȅ��L��/&<�\��ܥ��n��Mŕ�PYG�EAg`�@7��爻XR׬�.�˟���j�e1�~�YQ��=��-�m�r/9=#�C/�,/W�GAF̾�ξ�ƍCSZ�� �m�*_���T�{5�l��UF_��Ipz��2��#-
�x(��C���/2�7@���㾫���=b\/A1NX�?�3�_i��{�K	r*�OI�5�l�Vͧ��nB.&��{7
�?qڑ���n7�ds�B �Y^�IVK�9�r(y�I�֪��`g|\�Ι��~{E��~R)���f����P�C���^�N���h�<�g�R���1�3qFz�SN�X|Ŭ��:�tS��-ɿϒw� �k Wȝi�V���t���0ǃm
��Y���j@�u���a�����ߣ�[�l8�h����R;i}y�e��	xU9R;�r�ҿ��a��S�M)��ə~��L�e��� ����/�rʃu�"z�Ҷ�i��\�5�O�jN^�s��;�Gj�Iе*2����|P��0�Ѧ���؜̠ ~l��t��b�K�wz�FGv�।ȧ��a��!L�K;�AF�>Z�|���θ��~�ؗż�I��(0h��#�Z�@It��/�|��.|��$Yg���0��}y(�T�m"Qq��s���<������������&�9�YȌλoj��N�T���s;ʴB�1N���o�`�9�M�a9%�(���D*�Ę�������c)��}�������+��G��{�f��+�Rb?���
h�u�R��d.�p������fb�O)(�W��Q��O/B߲�k������>o���라��@1���0;��SFI?Զ����,l�SLgve�����'���i�����$��s��XmY��y2�"�?6��������}�����~�:|woB���R���/Q�%4$u$���A�E���N
�"���1w��Fa+Ӄ���Iױx���o���C�5?tVd�q/*�s׮�<�,Y�z<[�חb�o��UWى�a�~�iX^r�H�����Gd��G� r���$�V����X�Mm2�̦�+K�u��~��W�_8� �v}	]Ǿ9����fT�}F ��w�/^ğ[�3?����>/��uec*u|�:|/���í�:-��'�K������zڂB�v�i��<��b��/��j� 7[�i��g81�.Yn�PőV\M���8X#���_�a_�ީ��ҌQ����ǜB��䅖��y���0�.�l4$5e 4F��,!�۳�_�P47��#��GBk�LK����gc���,\o�w\�`� n�&�S�ߖ�|E�Z���0~��^ܵ7�:M.����2��7@���<�����<L���f4�Ջ�T�W �����G�Yz�|g�Sd���s��,7s8��0>�Q�D���p���PJ";�0��T�K��Dͪ���)t<�Vߣ�/��>�NT�e@�� �ì}˲��ƥ}z�5`��2�{��*�)$/�ć�l�o�;��F]��M�;r�M��>�@p�LZ� �q�EaW�u�s�F�c�=�$OI�q�B���'Y�̧8%?���4@ʞ���+�u������O�<(��|u�J����B�
�{Yu�l:Ԯ��oȄ�(m�.pu0<�\IU�?�j�����\B!����*�{��3峘��RcH�����b�����vu6�Q�h�C�͟Ø��6[���+�V� ��/�]�.��FG���Z9TCiF?k����Zo��t���Y[|���$V�����SD�i��c^Q3_giI�,{�8�1R�4�: jxg��q#�5?t:nz�F��;��a,,+������J���g �@�F��Ђ�w���|V��q:��钥1��Tߴ3��˳|� 19�*[��|V��8Z����o:�H%�<�j�.M_ԫ��"����KP�d�^I���-Jw�ˤxd���!���E�����s������]aj��:-E�c����{y⻃����ݬM�I�;�i�ڗ����Gv�Pgz�0��2��?o���Nvʀa<%[%?���-�RK��)�W;�����1(��m�X}��8jL�&����}�7��Ӝ�6:ż��� !;�&�hjL_����KT4;�5.<9���x`˞��rݛt���e�����r/0	iS��1���6z,6���^��[YÝ����D�P�}̋�p� �NQ��Y�f�T�����4��-O^�P���gi��Fb��nE���1$$��/��7���c��8k�֨��]0SecJMB�(�ڮz�F� fH����!�=�I�w��[����0�;���19W��C�:Xi���A�0��gSU�"�=x y�g�^)4'ow(I)G/�4�D���)�h�40���%��X��ֆ��EN�bL��^&����R��L&���+ .��i�ϮS�Nǟ3�%]��J2n"SV�W�e��T����8�%['ҿ��@�ֱ�����D^u�x��#��Oh�����S��ڻ�Gh���*�J����o���q��6z+�P+N<�և�N���3�>!�N8�:���.hQ"c�C˱)��8wd���N9�LeW�{>Cj'�%O6�T�����e|�_��	��S��H��⹓�N>�ҍ��0];�i�v�3��S?��]*���	K!�ц�������_߀��x�^#Ѧ�|$֖y1̄F�!Cs�	�u$ޔ^5���$ldH�o�R�u�s*L�5���%�Q�*�0�L��'*,'�3w���H��K3!���$�;&Ի7�z'¥3�?u�Mvrs����$-���!��.�Q{�"d����0�̢.g�(��	l}����A��uy��#��]5���C蝸�|9�Ѷ�*`��=�Uӛ�1���aeU�P�v�7q�K?ǘ&��m�+���� 7�x$�|��a�uS�g�%�k��Grp�#���\������_9C.�R�O��Tp`媡�m�n���k-{��*fh#�h�7�k�����Fx��uw��琯�R\�rDaE8�X��}!!l2����^����bϡ�Y�VvlB)��i��b�~	t��@�C�7p0����@&��]H
�𹒲���FG%拷-��wʘ���cZ��̂�ޜ �|'�'��i��&�H��K�j�d�(x�9�Ҙ&�T8H�4��h*�!�W��ޕ�C�ݠ��]�1�˛z|�OD��8ͮ�_���D1��L��
41�Q ����Ķ�eJ����//���U��G�$��$l�8�y�(S��9���*���j�ݑ
�m��C�+���Z�9>?��`��ɛߚ�� ��&#�.1�g1/�T�i�z�Jqw_wflBeS��sb ��*LT[8�$)�Њ��� "@��]ꯏu�9��&�D�F᝽'!i,�k�2�Gn�w4E�E���w�#cv9�(�H3p
b�,Ns�7�o*�j�r�_��e1_�E��YGG<���vN�9�z¢ג̂�YG��_h�#c�Z�⃯#��zQ�n��m>ַc�oVY�W���J�jƹT�`�	h��IM��9�ڃ�[�w��8�FV�̇�9�'���4�:J�B��_Ufu��sOE|���Z������g�e-�0� �]�J���Tv�Ghu�#貤�X�d� ���U�)���a��&F&�jؽ�P8/q�����˾��x�2=��I&��
��SԨ#�R� (f�m	�eEӕ�h-0z�(�YhŦ�3���m�����^��{Z�81�n�2�v���ԉ����E�T��p+�4V�]Eybyb5���Oׄ����"�}ܦ��,%#�S���!q��6u�Bj6]�-���'#Γ�4��.hiXl(�SJ�S��6k۟eo��a½ `��R����4��rKN��hnw+w����@H�jNw�X[ֹ�U����|QV3�A�R���+�ގh0d�Ħ�i⨙�9~��W�,ރW|�|��'��z����0�Dcڴ+�p��GXG� �*Ř�E��� �+�(���'t(�^x -���ɻ��l1W��RP�-Npv>����%�2[cp+�-D��)�4�у���x!
�c�~�3��d�,�U�Is3Ъǫ*�EÀ٭���" b���[��L�ʀ��Y�]���=4 �u��u��+��e۹�אj���l3�l�L(�0�������p�x�����p����U����%T%ld��q�8L�~~R'?p�����4��0��!�L=e����8���(������bn� M���<�:+AN�S�B����	��҉}��Մ��(W��.aO5+�z�GK�ie�׌�If]9/p�𽲚m����?�X��.z�� ��vq�ev��"�h2J
�t�����p> �*�k"�����|���#&�[�Џm�=I���]�K��0vj�.��2���JO�8�ś(sФkӧ�
��y�%�ITE�����J���'߱uD�T�/QY�+�<���̤ey�q���6 ����7ưԖ���r��$6F�q�RU��VjG\��g܆_���QQUN����>�4o%��l�*�δ�`��%(���8��!�u����w<'	����= ^�����a�;�2k}ZxSSC�����A��K���p3Y��ӆwxr5)2��}��A]3��P��R��4���"�t�2�^V�_ N�~���N�n�ҷg8��_�c�fR���;��#춋dWpE�����B-^�����������F����:-C��Γ��I����_q�	JE��}�p\ry�Qz��E&&0F��G���`rj�C��E�YF�b�-�v2�O�Z-��S����Z��2��v�����Db�^���Dz�ǝ4��ϟ��b#��3w���/(�2�)V$�������񂨡SZ��w��=()�e��$����&0��+�`8k�~����e����y�w����(�V ��k:� 3��8�l�ԓ=T��DV�iP�0��cM2֧��;C�q[��1����������z���w�3�J��r\��E��D/ڠ5��]�,*3��i襪!8 ķ%�_`�YA]ehu�"U1�f\��9&K�����7������dSU��Y;������o�Uk�^���V�Ȏ�N.�=�*����rr����d}9�L�3Q9PXD��8��q`��LB֠<�����l��!�}4Qn\����_l��0yxZ�`l�������H�/L�P7�����!ЭI�wF.ލ�����U���ƨw��3Й/)l�;ʜ}���#�xF��Ֆ�]���>�4v��OT~=�&��$Od6@�n� �BU�*�d���^��.@N�	��|
0 -�oq��j�)�3v����|.kҖD���6͝}����PЯ��-���<&�I�(�Y��~Z��;"f���ր}�,��@2���c�ZE�c����P��#�Dk���P�p�a�%x�^�U�J�F2QQ�m(�]��������#�̪X����?����D$����}(!����?�Q=|�,�	�m3�r���a��K��ml�Wj�Vi�݅��,�x�~�=�xg�.4���W���m|�>�`3!�F��F�fI���!� HP0�i	<A@�I�-5����ߴ�%�������h7`�������9�ʵyc������q�Bs�{%�"�-5-�e�키,�^KC[ɒ����T
�w\Ihk���B �ᮣ��$�ƕ����p4����=�
a\���g��=qê�YEb������ �MT'q
Uܳ�M�@�]�u��H���.X��z�~��:�T
g5�3���R�^nc�d��vrҸ�F\ǔ�p|ĸ���(;��2�ȹ���\~����p-�+7ST�=*0�߿�\.��8���F�|�'W�)�bF.s�Ͷ��f�˶��Y��Dro���7��7�l�W'�r�_�|��Ot�E��2q3K˨�`�S��~2�Z����e2�����dZ��^��9�gb���}e�_���ǜ��.Ut�r�7�C�2������8�-y�4��!�:Z�	�*[Oz7$/���e��Iv�|��v�����
���'c�(��EC��VJ��d�
{>�I�n�ڠ�X�T���V��Y^B���Ujxx�? �ܳb�W�Igj��׺M���}��'�/h�"U �j�-c�5g ��Œ�m�k��W;g^V�9jY�:TLm�����f8��tJ�$0�d���_e��i�ˣ�ۥ嶷2�b#u��n1�o�=LH2�Q���./u�iP�.CMC��k��U��
ٝ0t7`����	����w����o�C�.o�?��L`����Q�JL���w@zubE���.dM� ��������G�E���S���Ҍ��E}҉���׵)��O��H���2Q(ri6���4~��KºeԢM�<rі�ouR&## m��@G�U�B��a������ⅴs�s��h��9�T,�B$��ҊY�ब����H��w��XS�"�C��Y@�L���0&��D�&q�q���w���Fpy�1��3j-��=��`0�O�qH�B�=�*�B�i>�*O�k;�6r[�Q�v)ٖ�g-C�ӈ�m3���pG��yomL��쮳�S�k3�{�F[�*��@+��cg��!�ច#	A�\���$qu׹�I_������T�܈s��>՗H�رć�_PGtrj���"����8�٣��O��3|��2�D̽�x�*D&�?K�i8'?;�����?��a�
xI*|*��i-{�A܉c��E����k
�C��'�HW��=U�����HR�Y�i�}�h�C�;����$m0|�<�IX�q�vt����\��bv3�$�)�?�f]_\,5�k�R�Qv��a�J����5�?�のqA�ꉤ�	L��C��U�,�u,/p��_��S�%C�,Px�V�.n�������2IP���w������Q!:�-�`���y����Ɗ&Gn!��6�u�#3�%B鉎�M?��=�� ,��;)�T�k�,d��D�ڸrH	�<�|GNYj\��d4
ϹH��'��t�s��g1v����zf���ŋc`f�[�/b\�*���x���e&j��W�
�v2x7��kx� 6%���1uf:چ����inl�j!�)�֓u:�b���fe�=���C���+i�D�u�ʴذ�K�6V��^*�IF������B����2j��W;~�b~F���׊(h�{�5�C�3'�ݗ۹�8-�mU��En�ػE�(��8�� �o���2���bÊ�:@xъ��u�k�_��"�/��5���&�#�]?����_Ƅ_�̨1s��5*Nwu����`��)���+,�D���i���]�8��95��#�OӃ�? �\F�Cߘ�
[�� +J\�.����:!(��?;�I'|�N�[�ӅᷤZ��Ӷ_'��OQ%c�c�F!�V	&OB�0�
�..���2�`ڙ|(�#$��'��0rn��T0P@����EM��&ns��H�'�}Ҿ&�5훿��	���6OF&+
e����b�aR�����6m���ɧ��	=�R�>���_&g� :o�t������L�<Y�}�෋�A��ǏY��-g�7�8�p��æ�$Ű5>����5!H�
�w���0�������q[�?�h�)��ʐr �4כ�aq[�zC]�is��<��Z�΀?3KNz@8�����Ut+��6�ȣW���H�c�y.�t��~xV@j^�r�G��;�.k�4�IH��a�>�t�CYt��{5�7��D�{7�^��m%$�;��jP:��j\�D�r2Т��O��q�
�Q�@�w����-�=�<�;��h�p`hb/��AZ��=����/�m��L#��c)�����L�L-�ʱ����W�?�ɥ$�.�\��z���w=���'v0~E+��`�GJ
T���F$�6�>�kO���MN����3�g$��(�C�X��/�E�����G'��D���ۇ�f@:9վ���H�˒�V#1|��I(]^�Zp�o�d ����,9��A8X��{��/��u����@�1�$U��~N��o>^\ z�0�|s1C��ke�ë�$P����c$�U~�Lޅ�J����l�
1�Knd�*��~��Z9��V���^r�N�@蘌 �@��;G���q�������l����S΀?M����?�KN,���{�"+�7�+N�m�vB���Z�}a����|r;�Ur]F�wGs��i�6)D^
������`Ӫ�D�+�M��;_��m��j��f�8��3e���,���B��\��(B`�t%Lv[��Lͮ��ƽ�v���J�e%�hNs��n7�,�Ǡ&~hp�����bk�4;[d�hɹ�"�J���86. ަV�\��-��Q0��>h��&X�^��V' �[o@֝zGꤖmw��@���y:�,�g�Gbw��S�d��J$U�Ի߄�'����~.xQ�"���/�c)��p�)��'�g���=��^��<O�&*%P����Q.v��{dy��^L/���/$4�E�44u�8)��Z�uޓ��X����~Q2i7�߄��#�;H�Vl5����S���\���c��7��W��:f�m͒j�f{��oH��H�"���[F��ƫ����P�OEE>=Ƙ�28����z��k��v닶�X�)���=RY��	i,�1q����jQ���nLY�jB�>(f��;xQB��N�@b���+�}�7q�6��F������r�(�k��d8`��`��V��T��넍4�2�]���OQ��bWy��A��Jj�'��柮�O��sՀ�j	�����S�k\(
� ��7Hϻy�w��)PYUR�HVk��GT�����dZ[^���ly!����&�}%]��$o�E��B#�y�tZ�j���N�m5��xY�3��1�:��g�`�������p�c���ބ�%<��1@HvQ�=ُE�mEϝ3ʩ	��Nd�F�n�t!��h:��S�m�ӥ������y���h܌����Xܢ����>�����u���6������7jA��!İե����D���<��9�mNd}�p%�����������[  %;�Od�f���'֝��^���sU���E� �|Gq�i��
>QE��@a}�bz�.�)�\J��d�����.S�xC�����	�VO4%�"�y�h74^�W��R��rXⴛyq�£J�=�(>>o\Q�=[��>�{�Ar��'=>�������v���6򡬘��Q�Ϯ[����`���%Jȕ�� ��zg�����(�<�u�A�|�AB;7��Kw�v�j	��]e�s�Ji����5Y�-��3dx=!�[�A��g���Ey��q���K|s��r�q�U	`(��=F�@璋�,��v%&��AE����6�t�r7�,z���{�f!����/�sJ�F-E*6$L�f�.bc�ָz���L؂��sO�]-KA�ZN\��M�(۩�+2K����k��$�arR?qz�h&d
L����Mp�Ͷ�Fb�����4R�������/7�*�U���p~m0*�{b�Nq��R��e��'�#e��� �^��8�������e��;��R�z㽑�¾����:�i�&���$�'ޑv`p��bZ�!�E�򹐨Xf��v0�b�S������Y80���T-�1uA�͐2b�%���%�b�9���!�-�I�?��ڻ�]a�>ˎ)zc{
R���Ė���"���d'�3*vIv��o��"s���I���?�,16F'�K�-�<�p��;�f
���O��:�8F4��VO�d�q�"��}���È-����VD����g����y�j�j�L��[�a��@�_�p1�����/�E�Fv#��/�.����P�@��09��4GN6�:~��RÔ�|����E��&�Ǎx6��;[xl�e_��u8n�����Ʒ٢7+�����B�C�cY�����9���ȫ	P<�����Ygu,y ˭Gv�ۢ���[�G<�3+�4�u�vY<�ᓶ�ծD�\!��>��#i%�����U���>��4ی�{��x�[��7j�C�V6�_O�� ��E�;S?���6��l:*���Y�01͠{�Hk�{aʨ�^>���Ξ�{<��5�|h��&��R+Wn쵈Y{�I\.1��R��e��{??F������1YU��h��
����$ǽ�dј��g§��*��[�/��G��q�% � 6Q�ދ�6yk���aV_���wAxm�"�՘�����)�aʐ���Xy�'IvL$^%w���5G)6?-g�O�>���X�
�}����Ҫ��돟�/q�>�zql�,)��2�\Z���fc���Ej�K��=Oｩ
n�^�������0/��ϥņ�ig��4��L�?���"E ��{�"�v�e�zY�o��}�0�U�"�ġ���J Z�[k����sء��
��Cj�pu7@��?ށ~;	 �k�����`2z�
�ke�jC�0=vG<���>'p��,e�p�h�(��Ww5��#*CB�J��Ҕ���LB�|�L12@�X'��-�C}@��) ��&�I����y>�p�c�[И��BКw�e0ߕ$������)����O^���ڦ`��� �f#�PȷS�3^!�k�h�B�y����=���zÂ+�Zd��/��h��;(t�����ة������Ǿ3����Zw4g����t�~�_^ '�9=�ӏ���`E��N��K�t�����U�
<�����$<&Ǖ!�ߐ���ǅk�������᭽�L	�,"��{������P��%�v��Ǻ��о�ta��ʣc&�Fr eo�� ��2^� ��h-~��?m}�a���/����ى�G�o���#�ūq���n!,�31�4U>��� �I�'^&�`�P��a ��q)�ˬ�Y��UsԞ~ɑ�@��IL���QJH
dR�]�j�pϫb�<�t��h��y@s�l�T�� T+Q�
۹W^OV�c���C���opLBd3�J"ύ���%�#��ts���v���r�.;$9d_[[��v��u�B����L�z��7SCc�� |�>
��*�p��Hr6�Z�^��M-7�@p~�r�8�6-�s���ųu>�������"��a�`��C��09��*�z������l�Z��#
6�M~�����\��n���� 
�
bN��#R5 �����A�� L���LJ|�ü����!l��}��nYr$Ӏ��R�� z� @o��QH.�� �b�f�#z�HA��f���/z�v�6eW� b	3�˷c�i���j�l
��!�g'Ү[~ѫG��"d�EY�2I��� �Z��_K�W;���)?��H���<,}�[��FV��
#�4UX<l���@ [�;CI�z>�����P{Q��K�:O(�Bq���^����<�ٱ�^0A�Y�~&�lO�K�$������`�hd��	�>qv��@�&o��bĚ���J!��j¾@$�����⺫�fM�f'Qv����;�k��պ�2���Z�^$ֵ֤6���)��x"�#S�~\�(�B�H84o{�n��wr�?U��Y{����}���W~���di�Ɂs�O��T%FP�2S�� NJMǷ>�ne �[�o�Y+�nN���2�0h(H�᷌��<X �D~kw������Xl_�%�gF�ka3x��Л�.�٭&,����#�!�7�8��iG�z7���)\�� ����G��8����e�R�F�{�8�]ݕ���< �[�=�䵇?5�pI$\��N���_ʶ}k�JPZY�"G.POy�a,��9S1XzR0��TL|��[ץS;}��؁�� �d}h�QR:
\�{���@\�u���Dc��ʤ�9�~f�#�4Ջy�WU!x~F#�e�̏&�HbZkw讉�]e5jo�`��"���h.�Q���9�e4����<Z�$��p[�sTB�V�9�/S�|fB���L;}W�|��/56őXm�����4���V|�$�>�؅�,ܧ�5:��)�L:�Vb�Ka���w��#���'�JkW|0L����q�7���A�CQ['5������Oz�(�D\��Zɡ�ã,Q\��b�\s��]�ul�fW>��,�,��ؾ+�4�=��7�f�R��L���XW�}VO83��ٶ�����X��{�����!+���D�B�!���w���z"LI�J�1a!����ы�[����Z"�?{S��*�Y�Y��D���8�С4�LC�����j1�ۆ��m	���G���wB�'���?�B�j0����4����%�8'� -�(����Y{r?�JY)�y�NTpsZ���՟�)t�B����||R�ꄂ���� ]Z�۟ȼ����؞�Gln֣�jvf��Y$�q��q�8�L�z�� Q,��`�,a4K�����Ƨے�L̖����k���&�d�*E{�+o?�F��p#�$�R��t�ܖv���6�?����AC�k4�����D�Cy1���g�e�)��:��?[��R�*=u5 sV��&ɕ�I'�(�C/�1.G�f���2�	��´j	%5^��v	�1���l<;v�7P7�A�2�b@�� ��l ųn9�A:��aR)}�����C)��A��wI�ƴ>]��w5�q`*��v�3�;������"R�ܒ:z��j�F�W�C�V`�\Hy���TǕ���D��j����y0����ӗG����O��{�+�eyw���]��Q,�+���!� ���j������Q/���ChY�b'�g&�,�N����@�}��RQrHaˏ���������K�9lX]�\�:Ϡ��N/��l��#�`~aP�Qbe�<� O�nҠ�����cC���c�`��Fjt����Lkͮ�:s���H�j�{��Y��ޠ�tC+�+ ��+0��N.?�<�<��BI�`N���^�H��t��ڴH�@�;#���Cit.xU=�X� @���Pp��)�7����0u��-�S�=ꍜ�0��OƝ����C&,�a*�'������Cx�d0�n)A֘h86*8�	��	�s�q���c�1�%���3AsDʔ�8�jI�h96��pI�WN�o�X{���K5��N�N�UѺDp$�L���+�4��%�����l^ۗ�uz"��i�*e0�L�5��>#���G��C�f� �V�80w;2Ǉ#'�\;��������ҪN�z?���1��x�Mp�4�Η8�`�
����5��[�]�A4�_ۡ�>G���A_��N��ʩ�7
��-�P|�X�.ţ�>4&݂�k��K"�_获J��fL�ۍÕ]�j)K�`}�����P�ڂוy�D���0V��m1x����#6���ȝ�w\�.����廡�����-X'� T&Fֺ,�G�\�t��3V�Ȱ�w�ڭ�̂^�\������mvRR�-ǎ��N�zp��7j�F*����o#�(j�]XˢC��q��c����Ev�������yi;�E��|�'G�g�}���(ɹ��)�n�]7�8�P�P��|��ط^��V��5+x��Z ��8����L��{<H*����W��I0~8�p�&���ޢK�%[*�d#R�y-s輀a��A�͂J��;&^����8�d�HP6�BDZ=�K��R�[8�0�Yu,�#ۓ	w6��Z�r��jup%�i�q���W���宲s��B���ra}O¶vEZ���?Y��[���K��Q����u.��;!�I���\.������vr�d�
���ZE�\0g��r���x>���B�`&���k@*�ؾ���fc�H`�G_'I������E���A3�Եu�V#����`��0��;�3��d<~7��'JD<�V��4�v� �LK!E��vϿ��(��j�T��M�朗�PQ�zo"��WC�c$��8����oqsf�V��)��U�?G�O�cN��t��BS� �C4<�f�v�n���`��Ѷl� 8vHk���0yp-؋�g��X�	�Y��aM�SVM:]z
�ì���l����*ؙ @���>Ԑ��b��+B�����R�v150R5�f5��ɝ��]G��h�9�����^�ʧY���Őw�a�.�OiK��oCFb4l���g��^�_��U$�V4los������3Vޣ���/�����I9_�Pf&f�&�k�Jӿ��gϗ��h��JF�R��Q�@&v8?�P��~&�O�@2���-�֊��@UK}ւ�9�yU�x���y��lΒ���W��_��rA[�^���4E��,�:k���ҡT�,}�sQ[�!:�s�����7|yOS��2���"]�t㮫u��JIɂ��N ���T%=����\�C��
h�$g�Ոd+�}I��1IPZ=��5����:���}�`��.�����UiqO�W}1:�������F8�%�{��߀�8��jY���=�����9��ݻx������/�k�A�����R��!̎�潌F\J�1��.G�b'�ό関R;�ҍ�:~�7�Dgo�Y<���$�1H}��D\��_+6���j"����-$a�7u���BT�GA�`�2!z)88E��2� G8lom�16�������6Kn#�rr�=�mc��GKǫ ��0d�����tU��aސ�o速�܇����ޫ;	 J���,���8�+WR�o�L���=��U����`�=s�}8c�n��������-�&�\B%l���_o��$���}m��X0�^H$|C�
Im52���#�[�C�<f^�3�!hc�!��4�{�J�����4�U�q�`�N�LV3�����~&]�iT�-z��_��o$����<S~lj�/��^`UϠ�hֿ��r���ġG�Ԧ�b7چ�(���ʊ�L<K䋠4��)����|�	W���*�lUr;R/~���4rw �B�r������uk��O�tY��J��i�u��$�UU�sY=��>=ΰ3to�H���HiR���A���6���:�iL���C�.'ci����3BVyr�'G	���g	��8!y�V}��h��,�� \�w�F�+��Pfq���/�����Ω��A:�����eh�@n�ė�(�u{�����Rh`�|�k@;���z	;0����1[�'�q܏Z�y"�F��	sS��>�}��=��]�6���5����/Ǿc��3A�}N��Z��_q6���T�mNY�3�\��.�]� �Nڤu�rO��y��d���t|D���V~7�i���8��3��q��z�M㗕���<s�QHꬿ�&��ĐK��'?i.�V�ܪ�6�������b)�kU>����s?M��8`J ES���i�ȷ�ڈ�-���@�kw	&Z��>X"�Z��mXZԺmz��+����-�_&U��QE��*�>����.��
��M_�6�dO�}z��'��KE�^&���P��45]��ip6,�]\f��y���,Ѝ�`�"�+�?�Q?H�j~X,e�0��*�\��C"N��_�JBNv�Ȇ�c'
���C�Gѵ�)AQ�*���nL��-��wŦ��K{_���}��� ��t�ɯ6�<?���H$19����|-��"��:�n�IO`��D�>ȝJ!�+oY�g���'?=�4@`�Nk�1���gО�ذ�E���,�U��4t�4=��������)|�t�{Ĭ����Ez��ģ-.���|�k��q���pB̆���d�]g$�u��T�F1B�ɰ�9v��Ab�m8W<kr��:�	����[>��|�k�ەD�M���{n
�@R޴�村��h֗Z	���~;����S�@3qE��)��0\3�s{]���(�%�8��ˍ�,{]�V����4s/�tk1���J�����b�.sJ ��l�g�գ���������s9��ո�=N4���u��)(�� �Fһ7އ��A�KEJ�A1?e�� �i����d[Yװ�e,ٱ�f8��o���G5���$��"���(]��}s�ߒ%ST��獗^����o� �e�4�'�c�������f��>��Ti�:���!Q���v���KS�j�Z�1 �Z��~`+@��;(��w��_ACI�I�����)	.��?������kK���J#��a}��� �V6�!�ds�y��@���	�Ϝ=u����>�.���X���w�|��������l�k�E̹<�����F��w�!A�|����s"�!�I���ia�����f*�\~�ߗ�w.�Ѱ���T6���60�.M!�l�?Z�wl�]���*���9Ȱ EvV��K8Z4��NÑn�a__���~ڞۨ�h�ʫ�c�-�_d��@���%����I9��(��(��Vג4�e�G�j��Gmv��q��������d`�I�iV��|F�{)���,?%�2�Z8��P$�_�?�OZ�˥��#����i�'�iD��]]�K�x�J=E���ǹb��3s�"2�lF�5�9������?���
qv�'�G+�RWv���D�X����'��ih&� �Ɓ_��e��� ��eK���wp����{( ���oi�eP+¿Z'8x�V�J�o�}�[lgu��,ߔ2(�(%���C�n��8�5�)���
�}�����!Q�ϼ��㮀�6ߴ��<�����1q��m~�ƨ8[�X_��L��pi��>C@��w��#<%,��^F��m		@#�?M�qM��ق� �v�o�N'����a�H�C�I�����1�C	�J�X��R+�4`�Q�Ǫ��>u����@S\E���\���C�I��4�'�`����*Yf��2@� �9��u��4���k(&�'}�;×f�'ǠP�M(�T���ҝx8I���q���!���!e@V�qI�=��qR���"��	�7ku��wĎ��;�tFcq�d�F�lb�W�6����(u��Nu�y���N�ٚ�|BO��j��/�r�M�&����w23��I:!����Nr"�6F�Q�x�c��鑠�fN��,�~��ԯB�Ǘ��&����m~��lv0흩'���\��'�_!���qyxR�C��]��Y�e��IY$T�`
��{:�P��l`��Y�z���Uoo+�ߴPf�p\_(��T���$�M����n�\������-�*1��}� }�2��;e�ܛ �Ʊ�`^'6	7�i�SH�[��x@�M�a��u[k2�$�BR�[bC�v���m#{�U�1h�^�M�^4�������M7hf�#d
nq8W�c�wA���ʔ�ճ���u~]��G�'�c���5=���dU����n�R��8giRCd2�?LAK�|mݵ�:7x%�l�d���T.��\�Q�\`�CĞ9��s����mP��>��/������I�<2 {�Y7PG�#��
dA8rڷ��(56�����?�+Tc��w�V"3@x`�ߨ��|jV�݌�W�$��|��'-y�_N�:�3l(,K��pԺRk�]�g`����x��ޓ���p�	������l�	��0��ֿ�	o!O#��1��H&I�<�R�w�!�b������-g�!�����lu�2֕~��%JR�(��nϼ	�%��K[�~��o���k��E��T3v����޼��"�D� Ҁ6`�*�#�T��r&(�^���a���f7�@ vZӛ\�I�ݙ������7�|l2h7*�������W{�*b���aT4�o�LmG�
��f��m��S˒�G�:*�Jm$L^k��yk���H����S���@}Ȑ����|���'6-{�V��D��u�k�Lc���:�J� `�� �rE����O�k���Laֹ2��>�`�+�$�?ͻ�J����X��]F)�M�2��K�L���0��������@�0��f<�lnCk��p�S��~�$Xx��0�ͫ=�>�D���Ih�{;��}�u�u�/���W%�}swV�1��.��N'�k#[{�ˏͻb`�,�A~�*hqd��E���HJ�5I�ЉFm�v.":�bg�������gBb��Z�X���vݘ��@$�^B
�}.�y]��F�hA eQ���|�$�oʾ�C>}�Or�{�u~�HK2"Y��Q��1� ]��V�#KQ��7SƳw��t�����X���`bg��A�s�����/�>�Y�������3����/fgL=}Z���O�����Tv��"r9���/mX��?9ڰl�qj_*����{�!��Q��G�-W����T����� =a�j�-���^<�W
�̲��E-�gZ��r��]V2Ƙ����KꠀwbÃP��d;p�XK�>�rr9{OB.�^Z�X�ߏ4=+*�t����U�H������G����ݑ<}�`mM�bY�F��3.Vf�S��^'�\�����'&���'��H�<gf3]OU�Җ}.�[�� ��t���lu[~�2p������,G��/tC�4��=����u
d﯍b����'KC��3���g̸Ca�����CX���3_&�'n�1]]ke�ժg�
��]/�MS�(����0���:������.����;7\���h�����Q��8�W��%�GU�oN�s�'G'�݄�z'I��?�H�Z+�Ơ��fVDE��B�4���ܒK#a�RR��0�e�1a�D��B(�n����Q����z ���7-�U��ʠ�A�NM:��5�}��c���=��������v{�㗣�È�Ι�j��e�����V��+���c,�6@$µEE��'Y����W�x;��i�6|��.��+1z�NkZ��fӣ�#� �W�9oIu�;�D�oB��d2�=�=,��lc16�
��Ejk�!�-��D1����o��Y���{آ�L;���r�dˆ��:��
�nE��&����^H��i�0	����a[jꯪL�L_�a��rt~!h.�|�f��f\݊��>j�ch[eآndv�iJS�PEG�A�t V��@! �?�����1!姪�?u�[��� %X��O#�cr���n��Ǿ���UD�t޸lث�"�^�8�|3�X�mzP�<��P�BlԡH�����U��_��3�$�4��P��߻<�`u&�
o��B
qut�_��)3��u�x�^
;�_ޖ��?�G��b9�\a���6��,�Zm�1��eY}�g�X}�hZ+q(ضw�N��[�p���d����O�+J�X�wS$�$��#$��)1
���Qִ��ʗ����
ry"a=����|X�l�e��:���yuԝ1�yGB+B줾M�Di-8yΆ�S���=2� �y�]��d\z�n���ΰdP:	��\ÖU��� �N���S�d&ud߭��,�4�w
%�i7�hs �_Vt�Iz2�kйt�f�b�V4 #C�Z�����S������e�1Bd�x�Rn-�ʁ��IK�a�E�k�x3~;(0E$y�ǽ�O�C _���=�j�*�>��yi������)��@V>P�n�%�S�ꄓ3l�!�1�����S���/mIV/���P��ʄS������a�3 �?W*�[X��@{8xA+?�KB$֠�~H���a�A�*mQ��Ft�.ݖuRp���+�v��q�paD� {P˾n���N5�9%�
�e-�_^n)0���,��zN�{��7 �v��}�~��C1k�����-r]%W��ZƧ��<�?-,��>>���Y�&�`?�������w�5�dOI`̬���\�+jR��?��x>ˢ���է��=���$&z���pI�'�vCy�,+>0p���� �{�x��b���v����ٸ	1���l:�C� ^�vT�u[7�C��h�����EH�׌ �cr��x�:���$mH�R�5�8���.:J��4?sij�c��>J[n'�.�e�8�(UǢ�&��цe����_S��Ǽ0i�!�� S朓+�ǁ���=��lr�V���<�@�zn�#p��IUiN݃C�G��7�g��� 灪k���+�r��ʵ�)��u�����Ƅl�X,"�(UCmzv���^l�&6�6�%7?5��z`�������v�lZka�J-r���MJ�~1�;Z2 �	�̱-	oLo�����NoL%�!n:@��:~�T�F�$SqT��6 a�|��'�,<ye}�O���Ia+VXe�g��J!$����8!��oC�螥�8iX�07\��{�U/ݴ�ЪVbU���U/~q%]�T����g[�0+֞��Q >�8�qa=a���3�b��"7����STߖ�wQ���=�$��k�F���t�[��+��&�6i�0��B��2�t@+��*���QQs+Qc�hGrC��ǟ� N���2�o����jnVc��xlΑ��\z�������I�F�dq?)mH���]���7G�뀅[�_�u8<��w�&�ȿWP9^!R�g�䠝��qa�T$?�2D����[5�۫s
�����>�P��(���`�X@�����e%�戰�����Ox��b01w�9�V_�1��u�	�W��lbͼ8�D�r��⸈8�P��4b���\�X:�c>��~�p=�0f^)Bz�_ښ��\L"�f~��MnQ�E���n��C"�t�i㎗�b2��싖d���B�?��5d��Dp.�^�P�E�@49�j"hN�\mw=�H��\#�p����TH�K4��_�3A?���slz�j���K�SY��<���$ہ���`;-4�nm��T\��(��Y����Lj�2��2٬���z���I�vY|B�z��D��x�F�и�H���Ճ��|e:-Z�g�  9���8��D�y��qA��j
�\� ��JQ��5�P�i:L��QQ�y��<�
��م*MJ�s}a62�x�wmsxd�<
��È�:A��M{��y
M��LLjA�(m��2�$m)v8lʹ�K:��I�*5R�|m��e��X�on�;p����"=*خY˖�-� f���M	���֒������7:�o�SAa��+�wH�cT��6o���I$4E{�i�Ђ�Mtm�o�� D�
G�ض��#�\�῰�F�-�4�tB��{�+vS��E��^御�����S�y�L��=b�h�،��K�-�;����H3��:��n?p�.��̛������Tj8]����ʅ�4��b���:����0��̑�}L������,�H��{F����WH���A���^��}d��B��0\�sA�U�.ر�#΢Xo�����&������&��=QO/���t�c�T"�!z�:=���&nVZ��� N\�t'���8�����x|��*%�95�H�[���|a���n3���_i����;�6[[j��@�u�8�&�-�V�T�����B&����$���H�7��w��җ��:D�Ƴ�5B������r�,�P�f���t��Ͼ{��όS����M�H��M�!+��9��bW8�V##�Z�R\F+����0
�nm�β{�������Á����4� �p�Gjn�4�].p��=�R|���v}�j��h56�`L�'��k�9�q��������"-d�l4���41��p}4ּ�g)���=���2�`'�x�I�`��U�X%��U:*���e�B������Q�:G���:��������+v��������DU�(4�ĩ��㫠�t.�!������ ��WE�"��.�i|���$�.<�t�RBI�$ �~������n6s�݀���vJP��M����j�`I8ԧ�(���)w�����߀j�^�wy���Y	l�ђ|
�;1�-h��	튔���JQ�ʱ�{`yh�f�6I��1�4#a*gȲ�KA�yW�d��
*�BI��ё�H�����޽��ﯵh���M��°_�k9HT?}y(�0�a�2�*G|֥������.��	����N԰��Rd1����|�U��\{���xjAn� ��,�t�0	��@BL|������H۽4��0u����:�'w�ςJ6���9��u�c�����Y	Db�HPF���&��t ��1�,Ð�����uHs˴�[�3���X�o��8n+�J�M����yl���!nv�8�?D��v
^���?	)l�"W�=(�Fq�YF�y.�V9����eP-���
(fy�D��-u<rF꘴��Q�J����HXw���k$�!aZF�G���#��p��@M
57�~Tƅ��ܦ;�o�z	C�)���G�[}���'N[�p��|[���5���,ܖ�P��`��g�Wj�̌lEj�AmE�<+>�ăتdg���~���un�<�0�[y0W!G�������׽060q;%e�4L��o�h�T�*�S;�¾�i%؜��e���`���8���3�	BX's>���ϰ����,_��N-<A�L&9c�n�-e0����g�  �m�<3g�b���� ^��XT���[5(, 5ٮ(����Y4�o�� &�~�:j��<FOȐ*[]W��G�Y,T���u>Pt���UǬ߄c]�nhf^I�V���?��� ["��x/;��^L����]�FvT1��+]�ML�׆)��ݡs!�&����?j����,�N����ä�<�I��L�_>o�<��[��vz*ti(����+����&�%b�_���b�V���:X�"���E�����E�w\TY�0�Q��Rue�%x��%w
��u��h�Kɯ�'	e2��[�,rh�Ii���?��ʿ�Ǯ���Ƴ��Y����J.�s}��W4���M����z�`&b���}4�۰�8,z�lp44x���l��gD�T�`��dc�P��-�.��7m�<���C�>I�[U�k���X�u�et�d�(�) ܽ�t�YWcl�����������dF�ӏ{���OuT�����C��7���Xe3�OT�U�zz��Kv�j����u9�(�-[�*�V��ҕj�ú�gU,�/N��\�~�{X�t^Q�\��a�%5n��d��8�I���piu:1��σ��Qc�UO�K�Ϧ]$Lnr�2E��Y�@o}i!A%���U8�E�r���������K/�-$��V�F��	�_�R��r��������XVk���|�c������l�m�O���\?�o���Yh��#��pmd##�/W��j��
�C�.�> yh�֤{�fS0�R�K��.� #��w	+X��@��~.�sq��9�����@�R�O��I��������4{��cP�紮ጺ(d�r'_�	�v��1B̲p�w�
G���SP})}j��9|�3�� �&��@�ڳ[���M�f�~����%����o�AJ+�bP��CZ�CÅ��0,U/�为%_0���<��ޏ[��M_�h��FG�a���?��D	O���G��.��4&���+r/;7��_�"�<�m
��`į ��"(�?��˖ �Aϡ�i��j�Y^���V�*��fp�Y���KFS�Q�S'�_ɤ�OE��,����*^zF=�L/�ї �i�m.����H{\l�5. �W�2���-�c����i:ѫߪ�^q�J��c��o���pP����؝�V�ݽ0h�@8k@�肨���V��0��ܦ�?;���{�l�^#�l�*]�j���^�,!}��kv�zX[L�_�Pf�^⨔L�w���Pa7�����Q�i����S�m������x���D��)��A�~\��).ϖ�ߥB<h*օ�K���CT����\~�V�`�f���#b�d�AK�/��V,=|����s�Ү���󕲤�@�ط�\�M�^�9�8�2��n�q���PM��%z��q���q��
_��6!8e6���4��d먤-�gTm=#F�۴9�&�}=�F׍�)Z��10+�����gP��LS��ڶ4���3E���5W��E�Gu�e)<o̖]��;��q�/|0胂���!&���X����5���DLY�sV�T�Y���M�M6[&�7����q�,���'DOLv�_J�f돭r�
Y.{��3bvδ��YןF)�N�o�덫����}�(<����BzTę�lP�1_q��I�Oo��wn0�x�mn/����d�%�<
�cޯd�F�)�`r�w�G�_��',"9E�#�)��	��!��NSE�����OT��Z�6�A��ڎXp����>{��L�wD$�b�`C��T��]is!0�I}vűҭ���h~=����
��WS2��
Gqt�(1߈5���0�Jؔa��Xt[	���LL��}� ��PQ�V,� 2���e��i��� u�ǝޙ���Х���}0���,���:��z��r;^ŀ��WPj&G���Ao�\܌�f��9|{A=�:<kN72s�.�6�E��ύ	0���3�u�qd��(� �LI��{�#y��1a��#���#5�3�x����K;S������Xc�z���s��� *��`��X9�*C쪝�h�5��(8�u�:�T�	ܚ��t8֯Z����n+V�3������)�u��K�Mw�pi��|F�KV��d$F�j�������asL\�+`P�.Eg�^����S�:6.3��BU�%X�(ñ�,	z��HSTe���R����%��7Z�wH�<�x��Y�yFqw�k��5gc��b�q-�GU/��@��R�#â��9�c��py�tr����	�?��SH1��&��@���xA����uV�p���=����$)מ���$���Hk;�C�a��O���QS�:����z���]��/�X�C%38_`�T�1u^;��m�)�&�-��L�lls�M���b�w �.����8�167� ݑE�鴔յFӾ=��_Ac�	92�[�������OF�&� 00u�w�춫K��E�ՠ��tezVqH]T��@��!���7�f��D��u�P��@�u��⎂�}�f�UƝt�8	�v�!�;�x�p*4C֡�ڬ<PZ�d���\����V�7���4������-Йwyk��_ �׭��A��{�.H[T�n��(h��j(�c�k������[�U��^� �<B�T���iX���J��7���f�?�DH���:�,�j������֌�����XӿB��c���m(,�ZǱ�,��Ƀ����Q���\�x��Ӿ�O�~�6�l�k�*5�oNu����9�2,]�X���4�c�c�O�k���*"B�$,z��NY8���I�������S�h���>�-x��#�S`Ng��-�c����r�� ��;ej��1-
�܂䳠�|��@� ���+|�0�C�8��d�niX���Q��N!�8���7V  v�)����)�]4s�z�I��)o��X��f����\M����x��W��+ ���Z1��l� �n>Ө�Fn:����B���N�O6e7�\� �� �iS�bܖO�����i���T D�R��i{hd��7�1G�r_��Z7����w�֟V�bO�hAU'��'�&��-Юa�}/e�6/�?�Ϝ��C�Ys��O�9�R$?����CL��q�X���?�t���^�{ݮx��Ň��{M$R��RɶX-�0�d�e�=��_Nc����Y/�nfv>_��X'����s)����|p��ҟ�HD��P^ez�7��p1�x�8_aSVo7���k����"� ��(s 1!ʅt@&
Q>իR)F��6w����.b��������o�t�܇FPٵ#���q/Y���{|�-�B���䇙�.ek�R�,�� ��!�<]諲^�J��*I��\$x{�B�}{3�ϣ;�n��\����\m1��i�,��L�GRVY�U_��+�/yR='{Z�,����|���۽�;��6=�)�[>�h��\����ʿMT+�*��l2+5B\:��S<���&p���ϡ����S�0Tw�[?��E$��ҹn�^p�%(\}�gE�=R%"����i�ԜJ�t4��[s�a�e�ڮ�Nt���6�]��):%�St=�۱�)<�}�{����}�_ �b�+d},��=<����X,�»�=�^����#ܑ�0	5�0��R��%0+E_}0��W�.1�nu-��W`��u�?�$�� �4'��`�3���-��-�G��4�=>��H,�����dN)1IT���=O��<��{��.5"�:��[`�R��_i�y����-�)v��V�|Ac����#��4�ɯ\��ȏ��\-��X�7�Rx�W?���F�Mn�R��8���JD)�x���SX��J}��»HL"49j
�ݼe��rU�����I3���j��G���_�^�����Ÿlf-�a��*p�R}�qN�Q�W�K^;k��	M��l�J�Lq�A;/�	����o�L+o���`�$|ґk�|�/���x���zVi�U�S����;�"G�J�<��z+���h�4a?F��c�vm7����޽�>��8 �j��W���DY�{����gG��֏�a[!nZ,b���EWTb�ye����o�p0]�N���*"=@�<Sh�'��A!&d]��z���!8,�yW��W�EY~���xN�����J�H7��]8M�Y�j��_�"�S�sњ��Ӽ�[� 2�J��YZ�k|0�lN �5�)�%<�ѡ]�ص�G���t�2�p.���}��j=e��53�&@�B�O��+_�N��:)�`�
+`�"���y�g�	����i/b1u���"��w}{~ŁB���mo�\g�Y�8��B��!C�V�O~�2�;��q�a��`�j2JW��6�d���J��`Ki�3_�r`I�E�'^�*�u�Q+�^�TT�ih�<�g��W���7�6�1��rS�XyVI v���f�yUS���]�����P���|����߀��6�y�K��`]aO;z{�L�VmL��d��x���������(�PM���}�Dȼ�š�7���zQ���*������B��]�+���6��%|N^#$���g܀ig:�{]ڒd��[����Ѹ�s�Aw�v���<�mm:��	<ڪF�Z�*�{o������ǁ�ݿǱ�,��){mW �@R��o��xV	Q�}o;)��v��^�A]:DʠP�<�.�� D"�O��VU�� V�)��>k�8���B�ƴZ�]�mNW;�G��6,ȅej��)s�.~�'�6î�>��?j3�����u+i��P�ƚ4u�
�^BӒ��>��jM.�����s��I�FN w�2ܒ��}J����q/�.����/�����'@�p�a�;Z�=�/�tgQ+Z�]�}i�ǭ*8�h�U
��홙
�jwzl�c�0܅7����
��@��Q�`"�MQ�53�h��}�P_?�V_��g�r��`_·N���R��s�"丢�e���.�b!�@R`�N�ш({
��T�?�x�y	כ&J=��P,y*��v<Ӷ�!V��5G�	�MxC�̷F�dCj)���t�h-��j��VP-H�М8e�@du}���tE{�wt9�j~)����O!�|dM@�t�ɣ5�`߀��60Tdr ��w�+��^�C��0�r,޳�SySȍ4/'�!RĀ�;щL���<�,�\k�F�*J��і�\\�#--�P���&���N��G�C��T7,�h��8m�����K?"�d���������Ϡ��x�ZJ��n��
��������/?�������+��-�l2��f64X�n�P�i%3���E�K�U7UH�BzHO�tH���%�s�	A'�Z�	7���lQS�9����:J����D�¦��W��]t� �?3�����Rݡg�ؑ&MV4�N�|4��}�j>� Z�Z���Y7g�(�!��8���╒�ml�ѭ'�x�����՗i���$'1)�)E�Vai�Q����##$sj1ۻ0��M��ө�<ב���`�����@�z,bD1Ѧd�Ti�d��@1��R�0bx��w��R��
$r�+�&uOS��4�/7A���>c�G�j'��T��K�'�a�G�ͱ/��[�P7NI����s�skx��	b��Ȳ���������ۥC��+����	E`���엻ہ����3�49"?B�&.7lgc�2P(Rm�C$;E&�]_	c��	\�	�4K>%D	g�Qxf66�
���r�d����&�@y��-�:?�7��lz��7�ֹ���nxb��}%[����B�䙊u77��j���nyN�ѣ�%?s#�CY�ڿP�A�ܒ~�4�*EKx��d�*��d�3�ܲE���Mp���>���;��Z��F2R�T�[9$�cDF1I�~n:�Z��@Sm�yW��]FO *�q����H�^���&P��N4����MH�����3S���� %/0�$9#*p��y�	UR/�D�Gk���XiRH0�yؕۃzQ͇�K�ݨ���|�nQ��fvM7��4X.�� On�����@0�/�w;0� "*$��H.�c_ۮV_�"/�~�3]p�
���!	c�\�*&�����n���[��y�7�&�t%�+�	����>��M��V:j�mF�ʐ��Y;&D{� ��]X��G�hT�#����󮪻(�U!���Xc�˹?/z��HQ����,Gq���
?^&���������Ҝ�Ix�h�Y�?|����N����#�0�py&P僔��x��:>��!����{��DL��œ��b���P��w�Q��N�L7��D����P��ޥ9¡����C.�>j�^��'��%���#�3b:� ��.U�otu��
9z~g�����PU iD�.�8M���!�1'\(��J�nA$@�x���֓�s�D�+2�P�"v�ƖE� �;�߃@D�N������5o�	�ޗ Cj�*�N���N�N�G���kWC����9@\w[
��Ҋ�_���p��0J�#�𠙁�%�J��^�f������'Ojx��v �P���:$��W�h�~�:+b݌,����
K�_.\wN��M1+����a���״6��*<���\��r:�#j���F�ŋ"O�����k��ͦJ�ٗ_�';�=�'׮��g�Y�}�:1(��m�܀�p3�.����Q�]&���i0���u�2� ��
Ĕ&<�����o�k���˙�Nۥ�;��}��Jz�}���ީ��/g�!f�(MNr�8�����g���o��N�9"���A��׎�P��bQ�li[�0A���a!L�Ys
*�U�/�C0�f��̤zk��&�V�}���e�~H��C��"O����ԢӉ�S�xc|eMՍS>��҃��dJ]��ݺ�U��c�e'��豪�_�"v@UhIݷ�3	�P!(@W�"����bkčlQ!���.����28Tƒ*�G�ce!��#g��G�Z �@޳��%�S�&���`eޒB\��2��#FK�jg��l�Cl8�h�PE����<��yg	rktn�U�ppB�ǘ	�4�R�9�Jw�v�(h*�x�'�k��r���~I3��%�ڝeظ����C�8��� ��5ɵ ��-���g��xa���+�CgiJ�Iy���-��hd�����n�o������O� ���c)�.�6Z�<�	6�6��/8��4� 縴L�؉w�	a~]�xTG�vӔ7��A�S�sB1��G�;�3����sB�>��$z�xc�L���01�aj�1V�I��([�����,;�}.��g4�y-FR���B�Q�����@g�����b���hS!�ۜ]���CQ:�֎g=�\�ct��ߺ���c��T�UP`ÿ`p|��`���.2Y�Mix�ޱm��x�'\��/=͡���!It��"b���\T���z���1 ���P�GN�h�XM��<P�/ܤyBB$T�`Ϝ���;���J����L������=���4�r����X��59Zՠ��� Y!�`y����@{!D���sFɄm���[�-�lw
3�*kG�)��q�36o	#1
�կ����{����`_��Y��*�Kޓ��(1�N��iR�P�߻e�i�iqE���e��q/��"�_G��\U�<��Ýx�U�z�/,�h�d�������o�����L�D�wa
,"�g�qn3�"^ڱ���\c���~&v	i骄!z)��*S��
d�S�Z�.�7i����L���{dZ���d�7j�N�P�f3�޴���b�ꥳ������ÉL3����:�o���Fu�<짏B����2*]8��-�K��8����gi�tx�0u�xA�"�*�A�,v��@B �w/��`��W��k��p_��[���{���E���-�]&qM7ƜRR߿{�'Yp� �P�l���]L���=Q�����z1�ȉ!rs��(��t���X>�kt�B��η���~��"N�����6���P�Q�����%��O�����'tk��s�br�Ч'>%���ʽsZk��I���T���\*}�c2�	�-��=ur I1���>m�r9�{�����FN9�s�b�hS��U��6�`3�=�� `
�⨑�U�vVRC�G���R*����Y�fgYd�)�^:����I��(w����&@��?�a���1_����ʛ�BU*���,� ]&�v�{���������pGT���z;�>,@p�$k��V��n97���̓��7Ȍ�T�SQ�}���\V����V�����?zV[o�&�~�G�T%�-u
#�fl0�s��b�pj�#l�"�Q��i���Y��e���?��ɠ4ܱ���.ay�1'�J�)p�tP0O��/���~| ��B ����ϛ �9_�	�-��
O���nJ xx�+����@_�I��~�ީ����12�8z�:s������J����Ͷ51�F6vp�^9~�#_�O����^15 �_ՏhĞg�f3�ׁi��y���.��nǽRc/QZ�I�/ ����{�����]c���X����W@��Jnu��C�/*�\��EX_�2f,R��m/�_m��vx��5�ax�px�	�n��oKa�}�	O$����!I5����#�X�RDQ�/.��Xq
I��{�k%3�a�9���z�VǱ]/Q�N�Yf�<�B��%��m���DL	a�8��������]2-��ۆ�ՏA�ղu�a֞��;DQ�Ыq���ID�O��v��"�B�f ��s�/������P��x]�Ն�n�mT0κ�m�`�2�A���9u� ��SrI���w̞����⪛��m�wAD�s�TC�ě$��L����;R���G�ue��Vgs�koo#�e^!2�{��{"��Љ�6~���砟K�����G�]�)���}���B����d�ut��\ dNγ��[���u��(�F\����H\�Q����K�b�s7��<#Β�I�d��A�3ŗ�(=/ߌ�N�\�T^f��Z�*�DM)��.��H��c��	��.2�GYS�+���}�Q��DR�p�P	E�O�P��*�/����@a��YYY��ҠaJ�����Ҽz�b�ff��x�����ڧ�W�
��O0u[�?Ww��p�u��Q������a��� ��)�2��ϖ ��}���;S��y�7k�e���p<�$���E#�Pgc��-b�iꚅ���1\_y6*Ӊ��i��kS\"d�c�5����זA�������Q$�:�{#@@7����f)�]4ET�g�fq�B�fb���]�E[������R����Y�~-R������wV-�(Д���с_�È�h;�Qg1���\��@����!"�҄��%zy2��iӃ���J$�^�����ݗ��������}�XB�� �_=@pk�G+����K� ޭ�{V���l�eI��s�O� ��sZ���'+y)Ь�	��N顈�r�=e���<
�C�Ӎ�.]5!/Î���
U�#d��8�<�[� ���*o�,�q[$3��)@�_d�|�Y(rCd%���������y����-�5���r��Z):X���;%;����m����W�7�X��=��Z'v�s�0�bv�7� �bU�t�:��	�jY���rj�'/*VS�ʶ��)���"J��V�&	��	e�&�j��P�01�P��9|���I�H=�֦��2���s��W��Рk쏔�G�\��Y"{q��Ȳw�P���(��,<�pP�.�K�:��.��E2����	�� OVp�X�{NO�V8!V6d�쿣��� A������H�R��P�H�mzD�x��	�"���k��و���3z�{��?�1�0��ȎAd������ ���b�O�%���+�@yf����k|M��)h�a�f��t%���jIr��~�ٛzg��Ҭ���B�0���O�S"RT�g�R�ɐw*�W�>�0�by����eV�0�Y�0��r,��Sr���4�w�޼�L��&j<��M_��uL���ԛ��iϳ�+��Y���O'D����p8������z �]�P��ӴY���d6Nq��䠬ˀ�>��߿틤,�|NE�T���V����G&�n��;q���+�Dɻ�J��d�Y�*z�B�5Z�WM-��h��`숞{���ޫ؛�!˺J���<�r>����&*d���E���|N�,���T��T��<0y�Ʃ+�|��T�R��t��-�G��w�eU%���塌+��g�vUN�'0g�[V8U��e�IK�*q����<�p��j���C�F�D�[���YK�jRXס�I�'J��#JU�xr�9H��z��W�~a�#AR�����Эh�6�X��kѲ1)X�E��H��/A�1�8I��.�nH/��8)ɐ����)1r���~(�͵��S�jd^M���X�Π��x�U%�T��g%0:n�5�u���3����E�$P�p3�#ܔ��Z'µVbD��m�Ǒ�h��m����a6%. ��-��y�鸑����T3��n@ M�D�b���OJB��{ym��O,�DF S�J'Z�ƿ�fՄ�P��E"d� ���b��-�
̪��R�p)�j�Nׄ^u�X5U	N��!��4��指�0�e�SE;�h{"A���֜zn�#�� �ZLO 	�*���r�Tx�l�g�d�d9��F���R�XO���4(򀀌X��P���|�M�_J����)��D,6'�ZYV�bnp��Q�C�+�����9�P�6���S�ӑN�|�rP?Cs�_�./�u�X�����d�r-ry��E�_�Mf�b���1%~���r4���P\��,��n�HK#v�"�����Yפ��zo[��J�.�Y}�W��3O���R��,Y�g�l�5.i@}�z��ULh�b�	M�^hk��Xz��c��_"6�vȾbi�G���$2�*!J�������_�ԧ�T������i$��́�_}0ӳ���b�� ��~"[]��n�%Q��x��KE$B"�/عP^( �;,�|<���~SL%p��Ζ=���ÌHaԛS��F
�^����]���)��cCp sH��h�.�*6�jJذlW�����G��M�[���6m��駶�6Y]�*Hr�,��q -Yo�E@cV��?Q�����Ip1���[K-G�}^��W3,I&��~X?�e����X�7e�6�<{X��o������;b�KmE)Ja3�ʢF���G���p�B]���D�R�
�1	[�ߣ*nCFh�+�8x�N4�Η�0$��B�J)�ҝ~�~������ �pW�)C3�[���fn���M�B>���A�FH�a��쌇��AO�s���e�-�>��M+�0�NfsR��O��}��fok�7�� ��g,��Fd��E�M����O��y�s��䨘q�:��9��6'W��]�7�=�!���?�E���а}�O:��6k4;����tZ�YŰS+��d��a�q�a�
��y��%��l��H�mL���+HMUc"B:��Y�gw��h�����rDvy�Qz.i�D;������m��ވ-\K� .�[~y��,"��G1 ����u]+u��D�]hg����ͻ�!O*�	��[�p�����'����[s��H�H���J��g����S%�c�a�����w�-��7���$��z�?iw:��g�AXk��x0�[33K)_���Oxꖫ�ak��u�؟)�O=���S�4�(a��EYJ�PQ����9lD�U�o]�� ���BIf2|���0�=_���{�<�tB�H���>M�������t>e��d��e�,�g�sd�8��}s��C�t�G����P;�<�db�.��D�ۈ+ğ���O��`�&�б@Sl�'�~�<G��/��&���Z�)	/b5c� �Л�z��D"� �� mlc+���@yK��֜e?�g�YZH��PZ��R����.ف�V��a�&�.%���'�����}��F���ci̧�$p�<�����
a���uPẠ���v�� u�;��ߵ~y��[�G禟��W/y�x�\�c<$�V(��?����o6�א-�����I�]�`�f�I.�H���h1��Y�֩	Q�F��3�eXM4	�x�o�01&&s�<�.�b9_m��y����pǄ��+8�w�����G#W���;Үޮ������h��K�,�1CΔ�S1�jbN��yM0CC�X��H��i��]�{{�� ��g[���(�F[�i�Ga��*�͌]�yB��Ӕ+)a��g)X��3鲿a'�TS�L9���3��2=N�j^9Z/0̒'��c�v^��\6Q��ߖh`��b��x"�ˍt����5Q�� �A�dy.�(��JaSu�F��\^:y!��{ϋ�S?��_؟;y>�ryx�*cW!A8C��L��ڌi+Ӊ��4aJ�����KI}�m���S~��/��.������9$Py��_�\6>��k��,�W�Ψ��1(^�P���g:{V_ʯ�)�K��^~�"Q�u�!���y��c�-kŶj����߁%h�]�A>s��r�
5�gp(���ߤ�ﵓ?����9O���9|C�=�qT{q<z��C~ �3��z- s[T I�>:@&����E!X�JF���?]_TA�g��i��1�i��EoR�A���P Н��8���U��t�Ӌ}��b(���U\���?l���C�����t�L���.u4N&*�6a	�²����9����Iŭ�iH.l���7�(�����/����1 � \���N6�E��ޠ�ξc>����$ ����˽�8xf�-Ru&��-=���7ۯ.��-]�����(pZz��xΛm����/����^���&.7V��A�ZP��ژwǚ�B�q<ȃ�+�;�<<0�6 Z,���?��` �+���?�����@�<Z�����/Tu���;�~ۃ�J�K*R�baz� 6p���+'@�!RbJ�������#�����5���ǝ-*����?�e��+��'q�cb��f�"���U�$�']A��uh��bՌ����P�%H�Ϡ�ǘg�ςEg
Cڷ W���@��@p0��UC�i�3�u���NG�<�'��a�%�y�ᰪ�ে��`u�s�^]��҇7KOZ.�� �wg��I]��^:��2���<�U���𱰠[��P�
����6��td�y?0&!?!�f�tY�P�x%&$��m3����lwz��m�g�q��)���\P|�g� Ж�k@���E?��+MvD
1w�jF�)0.�_��B���$�R��׈dJ�n���Fp��7�('1��&����HO�����=�8+Nk��;��Tucb��n�^�TA@p{�a�L�Uo��4��TeX}pB��W�`��6�IIf��o�T�aJ6��ƚb_ZP;�����4I�%�=(��8�x�ִA�"3��)��<{�)��5���sr�S]��{}�9��!����\xOϬ���wi�SVq8ևĴL���0� ��IA���x[t��lD�@�Y-�͢+�B��(x��ٯ��7T�`�����
~'����J�r�����j�)�P)$���b��(�Tv;��?f�6�쵎�� G��I��b�Ӏ���b|)a]�wd��S����}\��'Y~�D��13����mE�Nw�;i�=���2'|��O.lS)Y0I������Ԁt�V��J�쪹wF�e(���7�ǈ�:W��ҥ�g3��tG���S:�Ճ��5�T��E/>M6���en�S4$�;-ܬ
�(?FǏ�:J��A���<7�5�EL`����_� $�S �k�w�*�A��|�RK����_$W�8	qC�l}p���J3�:�������� O��V��=��O��Bi(����6x�h:���1�.@���il�ax�b!���c�	W[����:�����e�g����Ȩ������tyS���}�@�Xv��z������?A˯��y^�J�̖ĹJ��y�)��,LP�|�U[�U�/���HsG��(2Jhˬl�ɟ&��t*�AZu�Aϻt��
��Y�M�$��Fy�ϧ`(Q��b�sU�ޜ�d��Q�"�|����K��s�0
YXˑ7�-F�׌�ʍ1RL�a�(H�%[����?�E�;����;+���B�s����wZ��Ϭ��p�_Et�X�2 (��
�:��uQ��0�z8O���k �x�G�U�}���q���$�CYp��sI��% ��]є�
�tI�������c��F>#����D:�>(��v=�s^�t�hmR��-������@�%0��e+(0���B�;���XYӳW���HS�qF�镦��2��Y��T�h��Es��.-��D 3������S�J�� �*�l�9f�o
��8��"�TV��t�y0�$�[��gn#���V`@%�Ԉ�$O53CP��ܭg�nc6������_	�u�(�߅��>�kgv#Z�~�Ǔ��d�%c��'	�9�+��3p��I�ZG-:���+N�77��,4�<,��ݝ�������,�	��﯈�����_%s��$�zq��K^�A�Y�n�*�����@{ܮc����#��뇻�Dq�~L�����SFΒ���~��}��9�-2���Azw�V��t$���#Ӟ	UuT���(-L�r�QN�;���K�/v�x�pQ�J����]���eY��la�¦�]��x�w��g�W<*
�m��(��ԡp�|��EnW�ũ�%���LX��j���q����.H��:]ب�9�UEV'�T?�4�B�:(j!�D�_3K��.��Eר���E������3�kՋ����I
�2� ��+b�B�K���&IPԖ�����]B2M|X�\�r]N����tM<.���*��fr�T��G���ظ�ϲ��FIM�����%n��v;��V]���g	�i[]Ѫ��P;�䧞r0'a�xG��8#j#��>�sj���w����/�]��<��^��<ݔ�(�����VR��s���R^��׻$5_�H�#5q�?_���'v�ߝ�!����*��j����Nu�R�>�r���|=�A%r�8���J�U��؈�Wd�ݶE���yv'���k%s���V�mے/�j"	�L�����+_�d܋��[�X���݇��הB�\��I*LΆ"ag߾!��$���:�׈)�nw�c�^�.���Km��d�{�eЄ	Q�6�r�J	�~�C��u����+�$���o�B� 
���I[c'C�������l\�_�)v��T^���"��A4�mx��w�(�Z�D�-�'H��-j��.�as�GS�޸WS:�����\���ͬc����p���q�˔F�gB���S�l� ��m2Z��8��_���$-Kb�bt�Ǜn��/�(�c����
+$ڦa��ՊıJ8�QS�ie�l�H�����EV
KA	�?&{�ҭ�4�a�"�WU2��'�U4�PG����K��X�rȧ�s����h+~#��ro�g5����D��Wv���SqI1#�ׯFp�reQ3;�?O|!@f%4��k��
*x5Í@h�13�x�[���o��� �)V����`�j��x�x�(�-�ߴ,�ا�<��d��Y��C��ddz
����O������e��{C����5���G��V�5!�{��} ��|��LL���#�,D~?�*�NT�����U����OJl7��	���6�P�Ь�Ƿ�R^
^���$z��Z�Wp6Vhؤ"������*x���G.�,��9b�xx�ľ"��j*�J�܀��ï>7g�Z��M,Kΰ:��"5]��`?��ԧ0�s��!F�G[Ӱ�N}6��6 @���=ˤi[hҚ�{���ia5Qc�@�zQ2�Ϡ�̡�9�[�s��m��{O���z77�^��?.!A�\��v���-
�Yb%�zG��}{���?>	�p�W�n����%AȦ�kZ�V^O~���^��:�kTz�=7P-gWzX�ɦ�(Z��뉓�֐����[>��:�o}@Ħ4ZW�J���
usX��K�i�cA0�"(]��؋����#ɗ<e�X��\&����@\y��`ʖ<�.
Ѱ���<�4��x޵�M֘*��Ls���_>bx��{"?���o��!i={l)r��T��P`�� �tUE�I��rx9-���=g���WU�j��R�~�a> �C�4��@�.^��(��΃e�	h���O����T��ϯg�Zg6h �V�	���+�/�J�Q���*�}���:�Bh��(g�F[hQ���M\��
�V�˔�:�ў�?\d���&�8hH3��E�p�����d����p�l�mF7RD�N����P��Iz!eC	���і��W�]`Y�oE�����E)Ӏk�m��F��ڜ��_v��\��8�ޮ[��B�@�i�S�q�dE�jH8A]��@�pZ�*Ƈ_����ı�"�Xa{5�ގsZF�"�e��0/���-5j��������?*y�ƛ<�=X�ЎJw�R��I�]x���Q_�ҽO��03,�+��˪�aHh�5F8�qA�ï�Ʈ8Zh� �����������7���)�Q<0��!��]L���t���(����8�L��1��\	3���jU�˹'��&���SV�z����U˝S?z�'p��^���2mk��Z�GpȇV���2�+�k뿡��i�	���M��
V�PzP�K1��g ����8�0
�&k��ɯC��I��[&m�5�u�Ji��#�~`�6
4����?a/3� �yr!i��%6�F
3��9k�`B=��VӮ�0.��ѫ,��`�� ���r�����Ν�+������6�q�*xd?�8V�&6�
�N�aEI�H� )I9�\Z��zM�TUrUˈN�v+�����}��0�sHЉ��8m]i�ڪD�(�.qm-O���F�.�@ĸ��?�J_�����}�^ٜ���s�*d��k�*h�\؇���=w�t�X&b�Zz�\�"r�E�L�������7�pD�rۗ�ݑ_
�i��5�<�k���q��V���2R?��n<z�X^/��03H���
%���$�(��]�@= �^lnD�%�Lo9�¿��fg�֩�>{$Bnwy�hYߡ,���R%�Z�؞Ge�ڼÿ���#�2���ћ�h.a⬢om�%����ڐ*\ryL�)y?��|�J�R��B�:���JמE3aS��32#�;K�n��E$j�qc����FH�UJ�����Mc�ƙ��X�TՂ�8��[��	ҌyR�'�]G" �6��&�!��[��B]vYy�b �g�qy{�@�zU,�ja��] ~=�m���ӡ��4��������
U��OC��T�=�D��������|�B���
�]�FQY���%�S������_a��<0*��ݓ@�ғ���qfe�j� ��x��WO���/������U�_��H6��b,y���͖<a�����%O}������<�|V~�l����{�k(��O��;Cf�o���vQQ�ٴpb�Dڝ��t�[z���p���ҹ�i�i;B$���*
S�7��OC�b;�tr�љ�ak�Fĺ�r����Vd�����
)>����X�7Jr��s�Q�_�H�@6�W�.��-���{ʷf�0�U.��'z0��I�C���a��lP�Ϛ��O�����zK�b7p�䳾��f��
	��q3&+��	Y ,��j��(�@`4w��
�u���5�7r�r���u㢠Y��G=i�1�\��P�"VN�D�������=˱���.a����`�F)X��9QI�����h�Bb�4U���?8 ��L�+�������a�V�?uB~?#�]����G��/�|���.��N�X���|�.�A_���o��R�k���k*��n�*)��}�k�l�m��7�3%����XB�؃��n�hl�z햴{���q�ɗb��M�	�B)2�b��\N��������ߣ*�"�o��GSC���(���@1�+w#E{�n�����(��������:Zҷ� �������dp��UC��g�i	9�	��0��@��^0p�Wd��n.9<��'6���R� �z����،wD嵍��]��gx��}���b]����qs�>e�U+�XR��f��}�Q��vy��y�b�3:#�����Ѧ�l�w�"����LBj�nvl�MB\F3��C����>�; �����
t�I�C�3�2͚`���5y�Dq��{᱊8�e\RB���˅�7�n�R���~oj�0�J��tlW:���Hީ��n��&�b�@7��Q�ҡLF��>�1��Jcy`�W�F����!~G6B���r?�R �Q�'������O��v�_��� 0����yf�������چ`ekЂ����߼9Y�,���4c[���*��aX�6������ڽL�� �#>eG%��գ�b����"����x �^�^�n�V��H~k��S�*���;j�e�?���i)�֌�H�Oڋ�����kⒶ�x��NZ�'+GY�h�T�k�������U����IM�jT������A�~��-{!��d�r�h�ta(qy�hp�_4Y�K (@�� �T	��X��q��ߕ*�تr�y����̫)�xh�\o�e2�L��e����-��]�3��&�y>����wYX��9�c�-�6<O��Dc�hn�����0^|_vA�R��[y�����6__�s���"C��bϲ���L,,qg
�g�+�:F=�y`!��z<w���8�ѱ�ȏ��Ҵ�No�Е_�n���?����iL�VqD��۱`��y�p3����dA�D���H��6\F��F~��dp:��nq���j��h���|�ϐũ;,F^	�G����i��A���mډ�:���h�S7��yZ�N���Ns8Q��􄧯��m/�A�k�:��8�-����c�X���ӧ����=�0ಧI���Gw�������.�G�/j�W�=��鿒>.�w�Y���(E�t0˳�T���"8:;���Թ֦�b�J�AUtf/�!�N�108�#�$?�d8�3�6���;h�O�Fy���!�i7�yޓ���	X�j0����=�>0P����+/�f[ 67���e�բo��֟�FV#ʚ~���$�򽄙\�f�4J%�y������\� �.�<����X��X޲��9�>�`�4��c�9�zm�~gS@��KJ_<%d6�MӌD�+,�C�����!�����Ǜ�ea_&�	0
����d�P��lD��+�x����^�;g& _<��j ]��I�-�T��-D]��'-�D8�N�O�Pzد��d~!�ab��ž~��6�-�G�4�&�p`1���	I�Y�ѡ���{��������E,�����TIx`D. ,���;Y�)6ߏm4%��[�A�N4���I�:�x�`"��(CC�[ۼN���t�R�2��Y�e(;�T�J��:ګ�����x�[a
��ڎܓ:����ԌE����r7��GG��?��as�F���J���hG�KZ4N%��B9 �&��i��%��1h��%l�� �	�֫~	�<s�����o�� �U��i���j~YR�jc"r.������K������x�v_�b�@ؑ�M��ͺA%�<Y@��bCV��쒛��6�2:��=�H��a{��G�c!�~�A)+2��F5��zu	Զ��r�'$���d��tv��W�y<߼�l���0��?�8BR6��;�y�yk�H	��闫A�,��<�~��>Q�*����Ә�R����^{��sx�"rBEP�逯0�y8 7Ƴ��� ڙ��4�"��m�u:ȕl���������m�';��s�5��@�����1�3��XM)kA'KKR� ��=�Ì��mG����C]p;C�?!���4���,��e�'�|���Z�g[��4���滼�gU��.16>���OB]%5�@)���x	��$��������({�n��wT��1ܤ����q�H��`oq,uV�%�`],�q�<�`f�c�A}::��b��d3���]��1�U��D?�J��M3b'IbFE&�"/�"�	�8x\f��-1�}��Y<V�f;zZ���E�Xɱ� �u�Ȥć�(�AR�b���~��l�Δ+�пvb,�5��J���-bk�b*jV\A0��l��;��J�DqI��t7:qs��t;�[�g���P�T.�̱+'���Jcp�쀽)$�'�(��))uy�E��]XTg?�Gmc%��ʻ�rK����Wn�
���H�UdD*_��=;�z�I��+Z(T��@ ��P��OZ���9�.j�I����6����9��f�i������,Z��ؼN'wP��K�Qt*�� *r�`z�H�d��i��τY����y�q�ďT�������68oH�x|Wm]��f]_V��]z��Bz"��Δ}K-l8wBK����M�Z����I��v˘|)���0B�u�Qj����qд9Lug#HM2_�f���1� �>��OJ�&�'Wk�W�tQ��NϚ4|b3P[�rN�?k�|�h��@��5�1:^)��+E�k��D�PW]Z_�=����Jkz�x�42ݍ�V��7թQ�6�{���xB�w��;��Sf������_�|P��$����T̙S�Z���l-�:ىs�@$�s�.���4cpneSvd�|�s�q��R�P}���=��s������Ix,�(����,*��;����ָ�x�.6]��i��ſ�,c�c����"����p�_HR�w���D�k���
�������#�k��	�ھr]n��֚e�ʁ5)�x�%ԁ�w�b�a�5���=K��m�#Tԁw�%/�[��e`ɟbj���g��XW� ���7.����������b�vu��n[�d�u�˥�1\���f	��<��R�>�ї�-D	��uX�U;����HU�n2���� O�ѐ�M	Ƒ�S�q5���]��j��%��rq6�n�,wK�p9�#�	M㷃胉Dt�.ȋ�����8~L:��t{q<���X�
#��U�{Q�r�§z�:�Z_��dE�P�T�8jEf�G ����(�Ս9H�|�'2�ºtkҸ��K|�x�T���P�[�l��[�2��n�m�ng�iϗ8Ho5����2��.���6qm�]��p˲�-��e��t�h '���Ž"7ӊ�x군>魖���Ppa�M��[L�V�
 ����o �|Ы�I4�����^Q�"y.qz� ��(�c�kbFф����<X�)l�X��|v���ǥwx��)���pY^��ཙg�$h�v��"'����,���^'A͋��� sv�V���������&�6x�u�	�-Z�t^��5�o��c���p���O�d��
!W������m�"���~�3�ű�E�F�߉���I ����F�$���Ȍ|J���ͨ6J����&W����~iR��ܓ��	�blr���7����IV#��=p���5]m}ׇ��-�ܼ槑v������&�ڪ��ӧj0t9l�r�f8���>�Gss� ��Y_��pG��d��}P���1��$z9��LK�
:��mq�^�'�NSjW�B����{�ß�?�n�M~�Q|n���I�?'���d=+fnH��]>�i�zo	���^�ծ٩H�_C,.y�"����P�lו���z�����I�*��?6�@��`��S���C�8aB��~7墏T��KM��?Ɨ,��#���|�/O�d-Z[O��yi\wbK�&�Mg��W�T$�Ec(������d�~����S�H�0j��"_<+8������!�*��up�M{s��x}Y�H� ++�0�T#����L��C����K��Z$��>��ߖ�99,A<�X�k3>�"q��j���X��QN��R
����(y!@�`�c�&rCz�.�fY���a���僘��x���k�p[����Y��k~��� � �������L��P�F ���Q��h��[K��L[��ݛ��I�e6��\1�M:ơ���.>���g(�� εj_��TvQ�� ����N�ag��,���I\�'��7�3a>�?�����t�	;�3�;a
�a��:q7����G]2�X�4�Il�PlK�=�%S���s�pBV��c�5ةJG"��6@7���}V��#8���A�i��cl4���}��]�伽[�H�BLEW��ٜ|�
�e�j�0��sz�F��
p������(��{�����K�]��g����n�W��Gx'���r�;�o�E�	 z����Eld]P8�ɽ�(I�i���V���������e�(dH�����*]��55�|�����_��[%��536��6��۞n>�?n�Hp�YY��G�AZo���>�$�2���t}�͵�פ)���O�O���Z���y[���y�U}�o��t?�V�<��������y<�2w��LesQ���L"!��LD��[O.��G��m�˿}^�0�f��/�!)@�ho�C�lɦ2��F�X"�fLM?���1��bZ��0/�?���u#J5����,�OE  �+���|0k�[�%�_����F��奖ڑZ&�cer�ڽ
��Q��֒K��8�0w�����@�.X,A��G,�E��߷>��#��?	6��(���F���6�\� ��OO吻Zy�u)���gIVsӋ��8�%�E�y!��ģ@.e�y��(�3E� �>��tĚ)+�g�MB�������:���I�����F.��ɓ8~*�X�Yi�܍�B�=,�"�W6��sx���k���_�@�".�hA�r�Q�xLLH�2�̽�(�����������b��gN7Y�f�),K&�%m��rȕ((x�U[�H��L�
��#�����_���{�TO�OWE���D�$�H�'�Gr�+V$�"cO���>��E:�Y|z�|��
��d##�x���$A�G?ރ���z&ht�\<wp�1�%�n"Ө7��$�:�Ji������1��,���
L�����F�1_={M�u��X�cN��#jp�0M��rO։ok+�j4
��w�jF~�o�������ŭ����"�𵲙w�R�'�+��8�!�Y�ሴ-���mmk����25#��I���"���_[�)�P�R��*6:5���c��1��f�1��nϧ�/C��Wmo�P��_�O�s���?��:��`/��G�y�!^�h&)]��[�?e���t�K z����d}�Cs�OC�{n���f>�-2)�c��]oI�S���Jp�Ц��{�mY٥:���6(���[1͝a4ooZ���}�Z��E���^.�� [������q�b�-���D�:����c�r���"X5y�+^���᫷'/N��迹j����ė�@��+�Vrk���f�~K��0$�X$y�/WE��e����r��Bj;Z�fgf��0��ض5(v���c3x�cT`(Կ4;$��$�/S2���-ER:�&6}�%o$>��@��E
aV������rE����k̼�?qp���SH�����߫�[<O�+ZX�k���奺�a�E����F��̹���1,���6�����j�M�;_��Ȳ�@$�������SZ��c*��
؛�M�q�?��D�<t� '�;E����Y:��4�Q�ơ����'_����z���k���IKT�*G�2E/�W-��ύ�&� NB�]F�mp�M�'�G|ձ��
f��5��	�e.��I$3��~�u͉����g��ej"���=��\ȘH���<P8��=���{$>Ӷ�ؖ<q�żAYɬ(w�
\�U� <�l�ݩ���M�>4f�h�+�?귔��T���~���M)��d��3���Bx����dc��JM[W�%Sם���Mϒl�儬D捛�S|���8��J�[u)k�|������o��ИUN�L_�u`�Ω�F��%	/kG�Wĕ������X�&f
BH�]�2@�!=�0���s���h�
��6.m��Y��c��% TRe9ceɛ>���ܤ�p��� H�kk>N0ĳ"�r[\n��&���I����9�!?F&{a�(	��n��%l��ѮsW�d�	�Σ�G�>����u~�U��e��İ�����������:"�!�'�S5�Ŵmg2ޭ=fKk��5l�̯{�lTulT�͖�xЦ��<�?�[�ŭ��o%�E���\�<3���:��-�>��c�MWFT�R՝���	yK��Ms�c|A��w���~���}�S�Қ3<FUg��H<-�xI1C�؞��2�=��� 턱�@��"K�K��k��!� ��]z����f�8=eʛ�1/�	(B�&����$�-���K�>b��޻�"�wZ;{��yw�D�z>gC��_o� @�c�Z�!�7i5���]�!�ju�����)s�'���j�CJ�r��V�k�
uݵ/���x3R�X��M��;��������B��4��Yȇ�P�ݽ���n��3�n��U��b5�/�6��=��)�<eWSz�"� l���l/?I&����䨢��S��]a%���K��1�8:f��,F�E"z){м?ZD��O�A.R�7�)tt?��S��������:{�_�ڳ:�'��0�U���"�~�¡��7'��.p�'���~y@�:.�^��6�=o����x�0���t"\�ü�iV�|�|�e���.�r7Q>=�P�� z�;>:����sg��NҙX@�w�� ��od�T.���q;Pp�L��H{���K={<`
�ocKn#�t����h9N�n�P]�}�����[��܀5?O�1+�P��&�@��%����D��m�I��ܢG�o�1�0��<�#^���U1@��R�qSS���C`]W�Q����>S����;Rm��h�!!�Y���{��B"�4.�4�Sz>t�fj0���{N��u0��/����� /�00F�u6yȷ<�՛D����_a��B���F��4�&/�\����Ǡ��I^����uv�5~E��p8B�V���Z���<��x�RN�Hٲ��յɴNu��ޟ�=���h�`<�����l@XӻR�RZU�]e��֖y���C�m�xB�!4�M��]��I�W
�p�ZǓ�L�qIx�K.=�F"�1mp<ۋ���ק٦]Moo�nk|��Fb(�h�}+3�E!So,HUdDW�w��	��<L[A�YD��M	�^\j5�ᚅ]rܷ�d'��D��0�Iժ@�4�2�߳��V��"� i�O�����̳���%sM"�X��]�Y�ZEV�qTie�
M��He{\|�1�]��=�wﬓ��6.�Y��'�6���8�2��v�Di�Q;�Ȋ��a�Z�>���bg��a3`�M�ed��-�&*7e�!����~N���wԶ�c,��fg�,��3L���㍯zwu�O�<���	�o���67�t<�AX�XKnXÜG����N�]>Y��z�ݪ�w}�{ZF���ҏ��J�9)�I٠e�i�Ā�ϥ�Ք0��O�45�k� ���I��jW�Ҡ��$�Ho�r�fD9��]Ai��ݩ9����n3aXm�ί5qX�@!���:l��yr�t,k��g��%EK~���6�=o��يC��B�4�O�&�ڢPQS��(�I��O��!
N���W}�V"�|K�b����c��"���\�����g�L\�T}������G�o^���u ԙ��hˤ�"�b"Vf�YA��V8���G�Ew�.n�8��(��x±c�l��jc;W���AhJҚ=9�|�blCu��P؃��M�1�k	np�aZ�v�{�9�cJ�)�us������ɂ2��[M+�B���y����"����ݏ@�tD�{)�������-�ρg>i��1
'�S� ���h6?��,����-owS�Y�iZ+j��p���*҃��K�M�5W�]r&��2���.���A
!%tu����ΑM�ƌ�#ť�nABp���`X���~=����e��!�%�c���Å7x�D�)�z�� �=R�0i��N���ٙ;HL��y6�뻭]���	��ZA���"����y�1�G�1�����isqŊ�
p(�ɟ�8C��P���1����5�lw��DX�R�:ҝF����╏�%J�;�@��l�U(V΁�e��)׍	�8����<q�L�tu�j%x0�N��r�ѭ�Q@�A�A��
:"�����Zl��������l����T���ʧu�Ȏ�Uq�N�`��KEx��Sl�#&�,�ܾ�x�7�����rԙ�eir��s�p������d�|����IR��w��K$�`14�L�,��~�v3_.�>rʊ4ϷM��2yU�j�  ѐ�3�@��[��-���|�Nyc6��n`}o�񢌑�ۉ�1��I�NaB$���Gĸ����T7��97�X���M U��NT�[�����j�1�����E�t��Y?������	<�n2+��tݕ�9�Yc^~~Z�E:qN�<\��R��c^�v*�St���I�)>?�� }H��p���̌�³v����˦��FǦ
��v/A75�Z�y�c6L�?!�-^k�,`��(%�ߗh��E��{o�&��ݒ5ޅ���6��������vȿE��-�kK�x��JC5��<%;lU˩�}���4h�܇vj�F���_3�V�%PkvJj�tNt��h�����_F��P��oV�*eՄ�3I�Z�z��+�j���yDEW�b��=�	<���S��$у$a�:�/-Y�ᎀ�����u��ϖy���M	1�zq��!Z���T\
�$N���'�����6S��1 �b"�@#��~�!��(b��8�u� ������U�F��e9-�*�݉L��=:ԁ�$����FN$�����Bpd�{�=�c�Dٕ�˃�n�|�Z)!rL����p� 2>�	:�X�Տ�UGzls/2�G�ZElFH��I���T?����[�����zux�lQ�3���6G��$M�ovu����H(@�}\�8w�f�^1?����~��=�V1H�D�Y���V"�������=��4+Hט΢\0�7AEU��y8#�����Ux;��*SdR#&`�Q���7W���W[�jSآN��F�8���<q���6��Z��uR'u�����m������k�����$���2;�]���.a��'5Ba�3��۽"�f+g�Wg�y�QW:��c1.SMS�q�f���Ν��+���2�9������A��D_����d.��;>$�m0T����	��1�U�~�ߧS�uh�Aɫ凯>�L	��F_8��%��OII��(��L1���X��"��yc�u���a.S�v:@�A�{�/�^ }��`��5��x	�{:����z�$ڡ����r3
�q'Z�ǜ��6�
@�ʌSk���8*�Qn��A��)����.}���yi�]đ��6}��Nr^Fʀr�Va-�\�ϩ���-N��ؚ3
��d� ;|W��UX����>M.��E��j�$������u�{2'kn���Fa�	r���L���6k3�_��N�{�W��F����y�g���n�:�s�Ly��BH�4y��,�f�^�u�����GchS������N��>����>CH�󁏏v�]��s����'��I���k%�v�6�~�������(}͟�`?>�U�5�2��,J\k`�Spտ9#̠w�ֈ�#�Jw�-0Y�� �ֻ�ƛRaٓ�/Sm����5�F]���)��`�d�3�B��'4�W�hFp5��4#/�����d"�%�\��C��Y
sh3�՝7�ý�����[ID��#'�p��B.���V|���^E�\��>PsA�$a9B�ӖC�kf_[�?���7��	���~�3Z�V�/�7P�R���}<ڒ��A�(=@�kj+�v�앝�x���n��飃Cn2��������s���}l��7c	�[+������^�PCϿJ����>��1��Ys~�7�G���%j�>+�`p�Ĉ�{1���j���W��o)i�3Ik�)�X��&k�`[a�i7����2�O������QHP?'�@�RkBK��Ak*&�q�>�C��Kt�߷���S�}{��IE�	p�B�㲄��us�R�����Ǩ�,��A�-�S�L֭o��hCy���e�l�	���8s�{�	U��1�P �|��>�8��������{�,��E�Y��yw	b5�-���z?b�x_�Y�c� ��~A�@�ծ�x���8�v*�ꄹ����bU��5�X�%6��2H�����yc�
uiuA�N���j&`���E�g��lU�[)!]ǵ�bm��]�����}d_�v��M�H�)��u�7�c�5'��H6;Mu�����*����5�@����GԠ�
mN1Q��ڊ��!m,b��_��D��G�P>̓���$�=o���wb'S�~cS=o�Ol�1�
K��C?Ut��:�8	���0�R�H���G)�mY��Jb�$�,�����dl�A�Լ��z���oKS)Ӌ�\޾���tf������C�"����B?[<�'�47��z�$�ԇ��`�p7-e��:��as��������)��ɞ�R�Yc�y�Eg3�~(aC��zē���D��F)��y�;A�F ntn18yQ��z��dՕ�
�����uW����J�a]�ۉ<Yi'ܭJ��I9c"i8�\�V���rF���F�̂>c�1�2�0����rk��-�K��*��a��=��Fc;�p�9Md�(k�����j�П<ݼ�g�AgA��Ý��G���MPz^�]�)f i#V�]c����n���!UB�����F����T;��>)�w��}��U��-�}UX�a��8��G���f/w4^Q�
چbJ4>�a����1!!%�K�l����w��ً��o�+^���d����O���u��\j�̓���V&�ϭ@�W��]
�{@��+vw��؝1RAso�-(8(��c�봺����?U#!�9�i��#R�2k»[��yݟ(ܡ򮏧rE���wN�
����`�'-�����Ʈ��*�[S���_�����$nj?��Cނ��F��A��'R�Z���ț�~��k�~�C��1RGj�ҍ:g�j��B��7�QX���yS�D���cJҥ��ĺ򭘱_q])(��i�<Ӹ�bj>#��<�Ԁ%a
k\��H���&rÑ�x�4��\Rm-��%l�|Bߊ��k�!���#5�+ghF�gh�@��j�HQU�4���� ^Q���T�lw�{�d/��"�,�<�؅-'Ƀ1iG0f�C����qv0���h��a��{$��3lc��|����tᾕ<J��ءpJ$�O-�;x�n�~�N<(s�)�����z����
��3P�g1^�Qz%�9���	֤L;d`��+�<�Y:~V���(Į�Sh�iG��c
f@�P�y��!��RN�	�m�8������2<���*�z*�#9�z��D��D�i���x_��uC��R1fȵ��}�x��o	���㏪ �ǻ���D>������'i�S�	���iֈ���2�=�V�Qg��q7���p�h�^UE�n|����^���񋗒!�!zW.9բ��3B?aO��W{
mn������h:c2?���DG4��|�u��}	)��_�t���)�� �t�^UN�[U
g�|� ����2�0��G���Ψ�Qnhp�fs-��	���O�v]�e�J���v���K���y�81=�W�b�_�5�&������)�[g���B�t\��(,a9��Y��d��Ռ�^��qN	W����(��_�=�W<5;��]�Vj�ˋ�d{U��n��B�(�{3�����S��Є}8"��a�Xuz����h����Ϻ0�� �y��:������̔c%^Ĵ�.�ʴ�5��J!/����"-�i_�����#q,:��rH�k��mԫ���^H��`Hse!���,��c��@��5|��z�%�g�1Ob˟�*��E�>6k�����z"hvS���'���:�B*� Y��7�P�Dk� ��x��A�Mʶ�8���[`����@�j�^z6�|3P����n�zuC�"�sߪ)S�p�#"$�lD�E�K����m(�:\V�}�Jh;m��/��X�}V+࣡+M6��j�(���	�]��;�{���T��fP�L�-WN�%~>Vs�Zψ�����S�N-^���7������e�f���S6��+� R[����^S^e6h�=�"<�f��u[:3�M�6#�}�u�w�K��un��$�΁�@Z�_���J�1�^O�1w�+��ڴ����Càx;�]��9�!����y��e|� (P��N}���@p�ޏ��q��£���ɍ��9���pu^���0�۬.C:�y�;���Q��*�3�u����v@bL��=�E{�W�o/�����}Zqp?0o�w�@�&��M����fB�� �|4��y�������w�4$�CF�,�e� k��5�U�����"e�ú��[E���3�$��|����oZ�\>ĺ����"Wn�C�e�7<��~��� l"���H��*!
�\�u����l��S��I�yx��&\W9+v�~l�m�\߫�.m���'�q�!"�-/.�I�\�e�[]%p�s$��0e��f0�=��i�D�(ƙ���Y���`���-uC�r?u�ך6��!r��e��3$���&8ɹjw�
Tj��J̒8T:w���m'!�_9�9��Ď-�}Yb�(x��_�,Y�`-)���|�D$tb2���)-��� �<(��.W���>&�����WEd��7u�D57i7,9�z��]Cߔm`�s���S2�$��@�	�vf�B+n�p�Ê���!U��������-:怈�U�H�4��P�9��I�]v�^��u\T�~�ǤяBhl'�R�����L�	����ړ����{]qR.;x���&ģy�ᔇmޖ(M�b�r�Vg�+�,�=�ӿy/�>x㟸����U�=WUI�nXF/�r���.�h���7̦2],]ky��!��ջ�@�W������.�V��V)��s�Ӫ="�,��?��Ыώu��3n���-����@$�����9p��ݸO�I�ջy�݉Kt��Z�h ��j�S��v��j/G��+���o��]xҳ�ϣ�'H�X���(�s&�S��eH�gNء;ڬ�b�h��4#VZs��/_� ������A��Tu^dj�&�)]°dǙ����� ��(0��餢�����(9gm${4.D��͍�_a�655'G����r2��*_��8
B�����K�qe�]{�!�UV>��7�3��-ReGb�Sݘ��[�L�1p6�Lb����?nQr�M�X@�
���yRܨ��Ĥ
��vcJ�i��S%װ�[{�u�m41�?��PKߧˣ(�����sL9ҡ������4Tl���(��P�3.`�i챭9~�%?]�Ş�xV1���r�˜�z)t��C�f�'���d����E��[���Y�e3���?3*(��EI�"�Gr�<.�M%+˟�2� ���c�IQ�C��W����I7���<d@�K��]g3C����^�"�'��	�F�'8������|�e�{�� �M#,�i@zʻF�iC�D�+)��J�;iW�����\|}���{C#�O��%�GK-�;�*���?��v3����7n��=�y���ĥ��p�f�[� �9�`.��{����gs�����:���9ّ#{&��0₡^�io?ELд��Fr�/�s���0w?L���>�]d+���gj�I�����l�� �I���"R@G
�z��a6�Ugb�5M�h��-v�'!����cŠis:�S~K����0� �4TgOS)��W ��qK���*�*�]����.I��'%��݁��� R9�m�A�pZ����&�Ӱ�GI�Ҍ�Dy*s^��^S�<����R�w�1;��#�����,�IhyMl�1-�	<�;!�\�˫' R:����Y�̙��-�ף;�MnzX3�ۦ�]��:�<v[�P���hoMt���/(5����Q����
��T|�U2r����B��<��������������u]���d '0m=>\�0���J]�zi��Y�5v��������L�{@�}r9g)��V{ii��%���	����^<j��L����y�Q�|
lņ�kL�j?3֏�>���s:��qa/A��\����ٌuD�]Ҏ�}DP�@ZW���9.��w�G6Yo�j���3����(�Psو��^�B$����H�Z�[��"����Bw��nLd��O�k���&��=Z���"c<�R�v�'�$<�d���
�b�C#�r�Y����Տ >w_�H�\Y{w�H���5-l<GĹ�?�Ϫ�<�����=7P���wX���݃��U?w��YPF>�8#��bj(�/���`�$��L�ջ��X�1唤�έ��#a3 y��҃ kL��ܱ\��מ�kT�k���T�:�وK��2�b�����2��*�4hж��cj��m_UÚ u���'��1�L�e�H�Ui���hk&P�p�fP7�R�E�H����Cxҥ-&�:J�_�.�'xv#�,��$K@ F�8��$�2h���' M�N��sZ�Ca|\��N��v���`�2E�C��l�T�7��O		Xoys�	S�Q4����Q�y��magm�`�q����l*��
hM���_�x�H��L#�+��^״����@��x�E����޲z6�RْEg��	��H1@���5�!���E@��P�F{��}�(�������_z���{�ss�B�@��v�����?j��:�80H�vc����8���}<Op\��ij�<�f���۔u�v8?/�VD�O��xA_�LrT�i���Xȳ�&�=�z.wXslX}p�����0N up���<0��]�����mv\d	Z� �!�qϱU}5n9���/^�K��u�l��UF%*�6s,�6|�#�C��}�y�Ce@-{��g)+�#`�0�|j}�#g(����mpa�a��#�A�K�4�f�Bq/_�[�r��@��-��/����E�� ���A1�]�W�:��ʁ�mT���n�vjun�o�:A�����W��Cj�jX^�%D��+N���C�0�|y];W//���]�A2�ŵt�ۣ�b��#�3��-$R��ٝ6	�J�vv+nL7gRt�c$��)�{vc��:�Jwj�j� �c1L�'Ӂy%\I����\���@p��J���Gި˖WS�#�P��B��ȸ�.#�5K��ǎ:���":t���?d@��{4O4r#����6�x1
�}4��H��j�cY�;���fN�.ePY+�[6i�M�� ���|���P�Tw��G}�7�Y���S��o4�Ġ{QOlFe@���H����]}�Ao)�8s)���:2�NBX���VT�H�[H�nP��B�8�K����z��299��J3躕m�s�a�5~������C�ր��Ua�v\8{�r@�� ��:���X�1cH8�v��0cCv�7��X�_�1 6Lw��~,��1^��:!`$z���`d�E����\�+~��%�&�����(a��l��Z8O�Ů�>6)��	����s�n���Kt����rH�V��� (���k� ]�).)Z��	Q؃x8W�e�I��$:���y�F���@�������U���i�����\'4�JL�9e18�3�Y�k�)�@x���/��Q��7D3䠾�r_���7k��k�[���>{��4��J��]X�_��yH�j��I��C�|�u3ɭ,Ư����,��3�qz�7'�6
��f�矝|�+��y��>��.��K^�{5xl*l��3d�����E]^��sNl��¡��̹kE��@""^�����tIL��y�/�u��_����Ȍ%)�w&�y��g��Κr�$�P  kW���)��C�����f��@���RCP|Wc��2)`>͊�ه\�X�"���ͪ�n0���8#$�q�R:[-}��o�����1�l̖U���%2��M"����e�͉7�M,PQC�H4�)��(�҉�x)� ��[Ƿ���"��`��S�/uA�=�HJá��` �����{I�z���gz�l�C�4�qD�����=M�;�׭�V���J���d��Ax�ب6O�8�k���Ԑ��O��yγG�w'X�����M���~S�q�oJ^d�"�^>�:H(P�h*JxP��w�C�q�
4���#A�& �t�f`�l���$����Y��%���/w|¥C]1e���r�N�4���XRx�S巃
����1`�����>v�u�q\͓�l
-��-����gڋ l�
�s�����R����-6\F_*<�������s֧%�$�
;��H̕�A\<��P���S&?�S"����I[��c*���/�T0�~�v�?���_LH����D
i������+Vj�c��5��D;���6l�Mg�[��b�%���v.���8\&(����]sh���F���,fA�L5���Gw|�)?4y�װ�r���(�4���� ����t�`������,�Ct��i��gܑU;܃��+Uc�$7�l	�ݦb���V\<�UW�@���;g����dv����L�%�b�u:/�ܡ�E"���y�_XqR;+i�&�
LL�D���w-s|4��!Z�|�"x�ߤ�a���i������g@��>|�mU����/����}�ё�H��_Z�%�uː�B�5�^k��<{_�nLy?�u0��5uJ-h���{���0O�!�o�TPB��mV��i?4�S��^ʆ˲Vjz�R�w�,x���Vo�≈���I�V�Ɓ�FLCC�tq�;�P��� WXZ�<��%�%:�?����	�{o@�;%[���oY���;A(0�)��K�'�`��	o䇵L�����,~��.��2���i�G՞Cl<��p�_OE|1S0�P��J-O,9-[H�H�C�R�'�s���(�����*>̯Ѷ�*fߌ��lІ����"�C�@���{u�A毩�Q���|��mAL�)!�
.�sp]��j��s�1��n���Kr�z._��Ô�k̔W㱎";�v �H����t��iLC g�՗E�"�5�ٮtn�����������^1��xz��'�?[%�nď�U�c�e��:Q�7�`QF�P�
�|�G��(ӛ|�|�r�H��R${*0#�2�T3�n"�ķ<\Ȃ+*@�FP�S��Хѵ��}�X�ǀ�Xp����*bv�J�0�	c�fRጎ۩�0��ܦ�D�~m�f���&�Z�{��L��S�	�#S�@��o�қ;b�F�!����fd�ۻ�w-P:u��0M_8���cy��g[%ˮ�v������{�nV��M�F0a�c����_�'?��A�x49��*���m�����Ys��'� ���0Oy�ضS�v���Š�
{O���R�I���I���q����Z������<�v+ ��4��������ٟB}k������>����@{�t�u�DU*?�.�?�x��M����r�k�SE2h�ʄ4%`��^m�12��FjyV�s'j%�$�|��V�|Vgi^�r��	!c��A�S|p�ب��b��X�8��^��}ܠ�v`7�RXx@�ɿ�����akb���ЁB,R6�5��U���EZ�8{���!������P���zl�B�}:�u�Z�@w��\\Q`����Gi,z.�r:(�z	�;�?2��ѸfRb	�7���? �bǎ�%���`�%��k��_�Dè��'�q���A)Q3ơ�d���KAO���N���zieR���Bq~����Ƿ��}��n�j�X�����q�V T�)����6�<���z��M����4y�V�vE[m��/��gs�t8d}��+O�Q��kXj�{��;��6�����j5f1ZL���=�_�4E�W��g�Ǝ��#O3��ā���Z|�J]���+��O;�f�z�ŝ��ky������ZB׵	Ь*��s�vg�����.�Fey*b��ↆ��K{b����O�74vZ���X>��5�d��cG��J�#sf�3���^*U��lż�?�vn-S�To�8�9�М{���C�l�s�\TK[s~�^�t���a�*N=��t�͢�7`������Zô^�|����/�B	"qd.iD����60��gA�ۑ�˲Bj�z�J�	�T�J�%�݇=`3=/1x\��Fs�oY�s>�p�;jW�.e��F�@��RB�e/���4C��l�
��H��w��Yg@_o[�#ف�Q(n�
�Rel��1-�eu�ʑk���rz�w���xa쁜��PJ��؃�dG�/�ʛH�D�O���+�1%L����΀<�S�C!#u`����6T~ˣ�MHNi�����}���b�yfy�<��(<�z���q>��5಻�J���^u��'t�����Q�A�ž��"y�!}_���)��lP�l�)��&I$����2�Qt��)�����t{_^�X����7�X/F��3vN_?��Gk�sP��DWh3�'��:}�x7�%�򾑎��		'��\�s��m��q�]9G���y��D}��z�H�w�1S�zp�3�"�`��?�G�B<"6�l'i����Xz��C��p�ö<�DH�N���rd7�AZ�A�Ӫ��	�*��g��w�@ݽ��������O r�,O�Z3�x,lL�v�ЀI*��Nk�B!擷�]�R� � ²�Yȓ���Ȋ��K<l $3Ǐ
΀�8��M��}D�%��W 2͐�k�UZ��> �Y�l۞Z���� ����2�~���1��U2X$<t�i2)ٌw�.U���o��f2���]]l���iY[����E��ji໋ժ��Ƅ��S���y����,��@ $=I��g@H9��$�ȳ�����W�]|T_��B���i��I��λqi7g_~j�෱�ޅ�zȲ�td���k�#�~h�J��)ɸ��ft���qU��Ck(v�_5��;���BdW�0$�����N13��F��=,�
� LBX�J/�R/���B/}Ҿﯷ���]M69�`�*�E@b�_��ɤ��z��K~sP	������+�o{C� +��s�((o���$Z��'lݟ�w��pŐ��nSX0�T�������.�8x�:/B�l�S��=�ԁl<x��x��桻ڀ#mG�� �u��_�g�W���߻KdC����� 6qԎ�LIu��%l"���
���$s�f|����#�D�'�p�U�4�є�c�E���ǽlo�S���~�_�PZ4i�����j�Z�c��W��������0�ю	�e�ب��T���;N�׵�qg��BX��!�Y0�����}�ʵo�} N�"m�������^�&5������ѵ���8G��0J08���ofyQ�@��s�k!�Fh$��TR��.�]�� U���p♆#"r��Ҫ�����:|}�jE�]8�n8�!>睋�����B~l/c������ ������:��<�l�4{�[g�J�����&��KX��50t>�v�w5�A9���E����芆��/P1J�v�b�G���2�sg����Z����%]L�M\��C��V�\��>w��p�
���8�+fM�k����^�`R���nm� �y�4`�)r	<�r��\�XY����f$��x%㯑�,p�]~m V����l���P�j�^/��Fc�߃�n�����$�b8�,�ʮ}I��@��z�	z�Xe?��+փe�z�5J��l�%f�ϓ#Ֆ�X6�ϥ����?�v�<q�,��;�5�j������=HVW��̓u�V\ʛ�$}�z�%�1����/&�Y4ܐS�����f�`&b���_���'\�_
�q0�3T��`e;��ʜEm��O���M���r3�E.���>&5Y��O�����_J��c�RV��.��C�J�v�=�=2ul�)�s$�6$yǯ�����.!`2���LP
�R��L�&��920>&'��[!թY�q>or�I�b�;V��˫n����<o���l��F(��v8n��m��X�����C�������p�n�bq�N.ڏь_o��Y����)w����K��W�iUI�bj�&���sĻ�e�ڹŦLզ�L���X��Dp�O]@G�����\S������|�s�+���Hx��a�g>�妚P������mL�E���~<��N-�*�$TS$����2f:z=��ķ6�A�-���U*���e㌥�]Zr؆��~N���\9���zl��r���d�4&d�pj������2���^4��4"��g�M�����Pֆ:���F�ݩ��B���V@4v��@C	�-"��%��p��cq� 傱}��7G2�9a�8|�ZqO�y�n|QnP��Y/�I�}��fz9e��?J;.�5��5���+��R���u���T׏��?�� �=R�|y�ߨg�D�5��őM���n[�P�*��*�%���D��o@���(R�!�T�'���?K���#����@n�YMdG�\��2���CS���~����{Tp ���H�4NDT�N�x�I��J��1V�M�d�$6X)+�A�VrM����,�r5շyx��Gz@c�ܡI]ń��RbM��3]xg�e�T��$����T|���9q*��Nٽe���r�B2��m�m.فn�(
I��|�W��R}��T%�7�5i�^_�"��'� ��9���%d�1>� ��#�a3^7Q<=�!/�4b�u�c����񦁌G=	���d�2<m*++�ŝ���4Xbc֍�)�A�q��3=�����s>�J�)��sc}M�p�	hBB8�p�9.Q	���>{�b)5'"����*�t�o�T;��{?%ЎPz �*:'G]�dZj�ת��n��Z;�h��>��3�r���3�V��k�N�=�����!�
)£�����4���b=���Q�;�����/�.���r�/@h	ӚS����5�C�lٱ�H����'[%�L��G���+9��4�
�|l�@	>e�F�II��9SG�<�q���B��S�ELk��Jz̥�����C!^U���19�^V�:`ܶ΁�CO���f�T��@�!�1�ɷ������Hap�?Һ�5�%�3�S?y��y7;���.&'��ua��p;���|�K�����/L��p��1kkdO�2T�P�|b�s��H~e���ޖzhR�����ț�Haٵy��p��N��1C���u]�ݨ��xӝ[���P���;��Jg�9��
.=@Kzv\�C��&���臵��y��Ŧ��eZO栥��;�+��Ɛ���pמŐ�o�5�� ����h���0�WqB{�7Y�u:����?�y���,;[��T��c9؃���0�j!�<�Q�9�,e�&�����ǿ�q�Ͻ ��:��r�Rt���eOX$�ƫ�{�B��� o�P^#���!G�x�&�	r�=��y,�7߇����^�"��s~�[��v��Hs!V��^�Uf�V�!$o��iT��i���5Q��*���?�:AQ�`#j�ړ����(I=F3�Q87z%ܥ,m+COD��a2)�w���S?�o2��BN-��68z�J5$�t ��95_�M��+�7TD�D ��vf:o}���=[�q
��Tr�B5�������"�~�-�*Z`�7�TD ��hD�|x[\��2q'"n���o_ZIK:�1��~~E�v���|9������t��a�YB�)�T�4x�QuǗ�����<�/D64���R6X��p�����3�=�P&/oc�M��y8��x 
��E�o1/wu�Nt�1	yl����X�����l+��������4OVM�́	F������VH�*������$��;;�3?kz�L�)�	��+"��
=R�����?�.��>�$n�H�l�q�b�5��T*�|�O$�,��Iɑ�Z
���0�+u?u�1�����:���^�I�h����������m��<��!1��F�*��k�E�vi����{3�)�B�4ۖ�K]E���gF{v4���v�
��>�A�<�}?����
��C�8�]�`����	P]���=Z2��rr#U@�� ��xPR��Iry���\�aS�9�Å�_���/��3�D�@�;��`��������Ze~���q��IY��.����v ��کۿ=��S�~?��+V�6�&:&�~|���'i=���ˤr� A�:J��ɀ��G"�]s���ٯ��N�|�yʯQby6j�!W����t��)=U,L�t:��SE�=tz]�q�E;�>�[�Yb.�Wg�<:9_B������%��l� F�x�:�	���2Ӯ5Y���\�}�� �`� Wc�I������\)K]:�p �����BrL��csQ9l|4�sIj��:�Π>�o2�<�Tb�>6���CNX�M$0��6�q�^�J���#�3�������gղ<վTo;-*�֓�e�<)��х�դ*�x�j���R�1D�/q�Za61�-��]���8�LD������M��5�����p~@8�,E�_$F��ݦ�� 7U���e��n�K{�K�*��g��+]a(v˗o�͎��ȏ�>�������gN%d��w��|����D�	�t�Ǌ�_a�߶�k���d�9��q3���"�@�yC�R(hP��������{��5�uC)|N�̮�/�<p�CT�ڏ�nO����8�+�3S�ښ2�j{,1�/"��B��NUVCbe%Ow��jKn�Y�Hzmfn�=�\����ɧ�"g܍mv71:/]��4MM]�&���c�K�PLg�qz���|�{���;xl�cK;'�΄�XK�2�OźU����I,q8����d����X�?����\�/�-[Ќ2�;޳�w{Q�
��:H������vI��L[�v䴾��� :�$�V��+�Gn�.�*0I�6���P�·�W�f�F^��ѵ���H���[3
�Mư�@6s�0���(\)���`!~��3^x��'���~a�串H����j�Ԃ+��9��"§�pݾ���̪.�)<�_�7�鑫������ؐ*g��Ycf�|ɫ��4�Fb�P\Vn���}�8HJZ6g�߷z���^
 �z�!uL{��}������6�б柘Q���DN}�`ӄl)�e���'`�e�>.��m�"�� �x��D�A��6G
J�D˘,}�rQ
p�5D��&� �a�������N!h;�U��.{>J�>m�7�dn{'�e��~�r>�xA�(5��K�$Θ�}��(p�|�G'<�k%��z�'͘?4֋����n�CE�d���OUZ�̓��wj�W9$�s��+.	Ò�3��ch�gT�Z��@�&��g��0v�oʲDZ�89�3c$k����&f��ݓ�AR�Z7Zl���-�N<��c	�{!��INX�ֺ�wN?i�O����6�0�Z�%S5�Tv�����X'�{�M:�٢�S��ߕ&M)�J�8�KÏy� Q&��G��x�y��D�"�3�Y�3�E��%��b�Ps�{P�ӳ��K�SV"�_j3s9]�b_P�T�'>$��S�j����ۈjc*�g��#2�����n"�+��h}|�����nf����{8M!/�K��c���
۞�/�Xէ1���َ%�H@~
���􍵡�>$98D�v��H��
�[�גe���eu$�ѧ񹟞I�S�%���xh+���A�,�+��h[�hz^�6/$���(�=�X#�h�65�<�9�4�8�Bm�Y��mE���kU#`s��,?G�9.sOأ]N�r_���OYs�:��A�D�q$�� NI$�}�$�չL�A���n�9Sj�[h��|�`����e\�4i�{�0|��e�$S��Wه<#�x�������M�<�`�O �����[�?��;��&��	��Tѵ��K�0'8��J��!^^ϯ�Q��P�q�����'?ة5�#\�"|O�Ė}�����+2���U[���� �n4&L�HT�$bnn�$��Q������}�%8S�u�k7��춐k�G1�W(IV�2X�9�>�pP�7j�,�E<��O)��e��rܘ��#���\k�&TфTv��<,�]9[(�u*C
��~��$��"����Q�Hc��1��A�Pw�9�$%��f�y��\5�َ��-k4��\i����.L ��4k�,9z:��RH�`�ߎgp�n�����^����f�qE:�>����#�8����#)�Cw��+�tW�9}M�������lB!��~���m)��6j>g�c')��=<߀C�Ak
�Lu�$�|k}7��)I�9̷#��m���LD����z9��:/�O(��BjgM�^�BN7�?���=S��b��F��*_Ɂ��Qy����c�n��Hm�j�%�q�����K���`�is��m'�n0���W|����o^Buݛ�% ��GS��S'����(����y���`8�S�#R��@��>Bw�r35��h7U~��Pf�˗�I��-�!��m��#ЅC��P�@���"('O%L@:]�sxZ(���I_���9Ѩ�֢2�#�!�cuX���hsp�Ӏ�JsM�3O؄V*�[-t1�0�l���}�����-6k�?�nK��n�tR�������V$�5mߑY %��Uh���Cwk�����!`y��5E��jϜ��&5Ѿ��:�X��m?% �2%�������{�$��ߙn���醛���c��<'ܚ�1"y�f4ںv�"M˔�,����_[[���Yc]"��
O9��9�`r���c�r62m�0J]u�^�=L�sE�'Р��Ի$?Ͽ�g��U��`��Z3����X��W�v��Sw��a��;� ������D�hϡ���j����� -�pa��t�Z��IZ����O:e�����v����9g��Z5T�Z�p�� �Vg�Ow�U�wDT��T�*��Y��3LE��$S�Qˀ���s~)�p�T7��o� �>5|X��riFq�lCV2a£a }��{��s���O3.���q�J��h1�|z��E/ׁ�C�V���y��"�E]�a���
�| Jt���i�Gn�ؔ*��61�!�gZ]e���X��?|D���j�u����'�iE�_�g�d�C�p�Qy�+�@�������,v3�3(���㯏>���e�G���*��j��4E�dq��
��X�-��W�K���h���A�2�5�УQA���Z�*� �QO�y��H�!TI&���sc�u��V�A*��^��l?����"
B5�ߓb���*f#٤�Ԧ��%)v�$dD���;��Y��s=j��'_�$|�y�+Rn�bc�]M̰�t�,	R���[�v��׍�	`�(�D�}QL�(d`?����*��V���f�6�������R)� =�W�4kY9��lɭ�h�g�K�b��kR��jU�A�襆i�k�G���x|�
'�@{�D{sU�� 51؎�r[b����Y%M|Kzz�|�$��W��L�������M�x"q�@񗳪�7`r�~���ɠb�?�Rh˯ǽ������81�\����HH
��JN��gC�M@���8�h��e���,����+���<[͡��͓�O�b�G+���igےE�\3L�ӊ��jܮ�ҥ��a��@�Tڅ�լ�Ս#���;�nɿ�`��R|�.R�M��p6C�>P�J��
��ps�OfJb�qgf��Ҩ�J]��� E|�L��e�C��p���Ld�M#�^ 57�ӻڏ͓M]�P�jsYSȾ5R�9����5�`���ud�(0U�w������]ж��r�a�t%�H�Z �4��	�s6, K�7��y��Y[*�,F���6�{�/R�B�i��|v�;��Pݖ����Z_�>�� �}A�J���:9�-*�5���u�n|��3��7`G2-X��D����!Q��N���4%`j{D5�����N�6ٕ�\n��� v��Z�UM���ic�ґ~��� ��!P��(�_�����En���S~,�ͯ���(NJ�J�э�zV �$
^J�H����?z����C#���ˊ�<��S��imɖ˂3Y��5��SKA�{�w�x���ȿ\:cH"�M��4�v(6YL��*��,~�;������V]�y�C[0�qՄ������_P'�]3�Κ��ȆV�AD��߂a���8f���ǽ�'ED�h������L��_R��MJY��x�oG:\�����6����mv琌�������X̣)�d���G��C-��q����f�ݧ��7ez��1�vV/�㮁P,@�[j��,ƍ��d�Jw��ϔ�f}7v�d� �$�D%������dGi������Oyvd�10_��> ��R�p���'4�.�'�.���	��;����A˧�.�6�g�s��1�}򷼶�P����[	�e��·te5����d��a��a֓�C=Ţc6�PE��0w;�{Պ��܃E%�7�Y���Zv��UQ�`�
�E��H�Wb���,�9��PB����
�I����@�Gў%�8��U���/�̑��2J#�{�
��4�DP-$�:'��a���
�F� \��A���@R�~���#
dW[�>�wS!V;~!}Z�eXu���"پH}
k`95bXo�эt�7�|��)���ym�;߿6����P�r���D�S�@�Y�1�3��r�NC)����=|�:k$	<=�l�j?c����l�I~%��A�	bCi6:?�\�Bev���_[L�U�f�C�"+�1n�[Wִ*�>�ij����	�P�ǖ��q�K<�--�;��<����yt8n�U_;>b~���2��ޯ��\���II��a��NT U
�#�C���M@ ���	4M.l��ⴜ^��?�E�ܨ��W�z�N�Z�G�Hˉv�k��QU櫕��ɴ���誈*a��I�x�β�R�*��M�I��	1=?�T��-f2�.���0Z���ܩÎ��������nB�b���Q����=='�ưlq�?}m�`�2�w������e*n3�d��-�B{fn��wk�f�,���:.d~�D@�o�w���SEM!����↕��)��=�����%zc^(��wxV������ϯ���\dĐZ���^��$vrL�����d��nF�pǨ�R���UD/���ܕ���p�w����l�l�>�dk�鏓�z}0�����׻�8@��D�m�� p檠��Q@R�p�~��AtR�p,���Ā\��k���USS��IL8������AK�2ف[	����r4E��@����6� ��Gn��KIck/"�������8����Ȉ����
4~������i+g� �!���q������/��oE҈�������.��S�S]��YS�7{8� ��w������]� `��-1��VƘr _��ga��cDCt����cJ�k�����%���� )�mZ��%�2N�����݁�j�ؘ»�b��EX�n�/Cv4�>�􁭹f�w����oIޗaW�L�Vd\�B�~Sv��N�6�2:Z( ����ѫ�����3�ζ�;�F$��4��y�"x�2�N4��P=������t�&=�MEJ"֟U~.�#3�"��;�~_���0��Lw�m�,�r-p�st(;�������T~ݜ�N�BQJ�B��ؒ~o/��V1뽿[�+��𨰆� ��<F���"��&���L��Um��\-�L��E��''?:�v��g�K=s�U�{	ҝF�/ �	g���B;�	�^#}��Z3�o�+�!z���L�m�\w^��-;�̩��'gL��cm���%rG����+?������V�`ޡ��<&cx����(��p.q)a, ��� _E���P
)��������zN*���r�u��Id���3.a3��c v��C�sꛔzu��<K�s���5�����S��Z�no&g�~r��Jm�p��3�����تRk�"FkZY%;������F�hz�1�L�G�`�H"�#��F)���	GZ���:���xO�1kTN�os����{Ι/xJV"ܨ[+�*���A�Q��*�������v���u|r���~�="R��<���J �Rp�Pր@F`<4ݑ�1�M��=�֕x�Yv�Ӌ�~>���Vԛ���>��%K��T6���nx�����@�Ը���;�"!Eȴ�v���C�ݶ��������x�����T��5�&�9���\C�9 ���a7I�-JŸ���T$��/�qq�^�x�r�L���0l�r�v��dw���X�[����i5"o���V�@��J7#�8����!nT��κL�0Y	!��>m��F�o�aj��5A�/��ΛZ��R6�H�=ȐٓЯ�j:��[g�n6����c�O�*C��܌Q�"~V��A�� �~��5�߲�3��;6�u"9�1���$�	����ӿ���E�!د�	՟9PV�K;�����+;Ҷ1����E���@]�'�/T3@k� ���9����m8�d{�P��>���r���"��D`	��7�u��wWԷ�2{ɨ��?a���b���&��Y@����-/�M�_ⱏ��H|�nV����<�ͧ_��D��I:�aD�`�%x�a̴�����\~�v����K�l�釬k��Qu�ި�ZnC�;v���ヶf�I���L��8 {Ez�(���dFf1�K�pe���Bt�]����wq�&nGOV�/H�;��{�(�(	��>OdJw�,��ˆ,W���U��z�����X�JW�<���R�N����9��4��$s^��!捱�X �D�9���#1�9Y��0:00��~5��{��.Y��̅�e�1�[����{�c��J�^<n^�kӏq�ݹ.w�&B̊v�1��_�[6��x��O�R�F��p��X<l�=(K���*�&[g�Rq�����E)�d���T����]�$�7b��[��^�� L;�K?'��Kb�m9�X?	����6�ED8=�����ѣCq}Pw��n{�9^�n �bǍ0$a^PZ��l>��u�iy�����^gpT�6��T�-<�ul�|�b��u2���N�C����
��*M�����T�-hLB��V�f��\T��p�1���HD�a�D�.mˋ8m�������U����'A�b�'���g(���zw�%�K���Ii�b"S��m��:�V��P9(������<`V��>ʹGZY��P��<��	gv���VA��G�}��挟�� !�Ê�٣$(}��	w��kΕ5��b#�9�]?�Ք�������^��.�B��;.}���U_A t�u��:z}�e���y�4u�P'7_5�����Vd;KG��4}M{���E-�`���_gj񥓿I]Q|b ���
@ dHz*����"#����l;ϟ�?�}+�!����K/A�+(�*Ok��&�0�x�$������~�Sy5�j�a����}��L8��7Su��	ߙ��/�{��*ߑK	�����υ]:�k/��g�T�g��V�a7�Ӛb[DW�ͯ��Z��9�v��m�S��!�Q:l��ǿ�\��*#y����}C�rw�{���������IÑ_���Dw97�Tܢ�g�O�>AgR��Õn�3�75�*�QXL���	t��6k�8΁Y��GiJǱO�.�����X�����<�V*iL��n�Fq�Ɋ�O�'8A&Z����\�.l��xk���28�$�i�I��T�/�=z�����>�ߓ]���.:�#�8���)#8��[��G�] 8�]9z����!�\Ïշ��V�\����_"���e-��T񧪷rZ.�݌�1P"}8�f�	��˶?���R���+���O��j�����	�r�$X���[��?x���~[������3.�_���P��3�jS�`���BP�#�ְz�<���ܻ�J<u[��y�:
����FV���t"���Y���� o����j��d!vh�HHB؃�:7J��@�*r�<���
���3�,"��0�R����6���_��Ljx�u�����vۡ�-�B��h΢j���F��f��|]�K�=(��uѴ��@�ȏ�&����EU~"|\u���ݽnR�N��F�e���x��#�����iQL��!�mS�xSn)`��候\!���;�����e����-01' ��n�5M�6� (׺�㎚��95���M�E��V۠NA|�cl-�M��D��X�+[���t[�R[�1�wGGc�|V?��|a�e~����b���6�ؐ����2�Z�1��5я�4���զ96
�0j�"*���k*{����V�i�:)�ŋ�� E�)#K�A�h����83
�_cS3Z�r!�*��s���f,��~�2��Dq�9b�[�����w�j�C�v���R�3X��v������?� � � ���w�Eiv����o{8T�mbo7`H��07;�^�J���<Ym� �h���嵳pyˢ6��Q�(9�[�c���%�"�CBW��""'w�h�����A��G�Q'��&ܜ�X�z�o��RRɗh�"�S�Ѧ1��H�Q�� z���;$�l�Ƥ;������Nbg�(�R
���Sp�,r#�VkTC|���<��S&h���Z/�U�P�]���X�-�f��I]��n��ˈy��sk�O��Z�Ŝ5h�R$0��q�l�	�¡'�<ӌm˒�=;�D������乁�����Տ9��;h����ש���%>�;^&Xf'Wwp��/��vc��|0���b3��]5t�r�p- ���_�g���/�(D~iU��(G�S��U�Ĥ:y�n"���#��}a!��U�1жҾ�LD?�gO�6�n�/w����G��� c�0���/2�K�Y	��0l��9�δ���T��/�0�{�kg+=��À���ݘ!�m��U}	
O|+�u{!T�ו%�\�2��<�6���=㺘��=��o6�"|�L\��=/�d��sAJe?*�_m\+���1=��Ի�G��=�3&��Z]]���rS��h����@�?����Xo�����Gc�n��[������갞j�鰑�w����lb^~պ��DvJ���J��,��k���?	�
U_tB,g�EԷ���˒dĐ�5����;��Ur.e9R�EbP�e����֕�E��������;�C҉̒9QhG.��QI_N��_���������R#��/�:[�a2b���y���	��x��䘘A�l�R��HV�ݪ��;��J&K�3o�6Yc��h w>m͇�����le�ts'�V�k����@�m� Xo�`�)���J�tL��4�R�w> @����6^C~
���K��H�Ű��yo���aGH��Kr�������Sx��,��B߅N���E�dB3쵺���@���\a�G�*���{Nn�CYy̚���a�9>W*4?�9����t��{����tp>�Ά�x�q.8\��R��&"H�������!�f�Z>���͢;f�n�����᧝	q!�A���ʔA�� 澄��s�-w�����T��&G�b�l�d{jn%�iˍ�M�Q{�81u����{O��e�V��Gl��*��lS����pq\����>tZ�,#��+�����ZZ���N�3�)on�h�E2y�(�E؜V�I��o�B(��O`;.
S�R�tca��{K#I�8⫔�i�B�ɢ!�SD�;;�_v�^��4B|����)��J���Ա�g�7�p8~W�
���3�M��a��;�a�O[��Jk��\Q�I �'�D��3�tJ~�jsl�Oh���隬P����D�=������J�$�jR왟��L�=����.�uu�|٪5�~RҶKW[	��$�)��D��dn�p��5sq���4��%�^A"���{49��K�==����1������&�3vb�M�r�у��3H��M��d`yv�U�n�։ ��/���y�����Qk��"y�.ؔ��,��N���n��-w�|t�aC�C�����z�~-������:��P����7�Z�d]!^�A�A����q�<�y�9A�9c��Yڤ�GUD�]�n�7���YF��\��2(�^��3\0zx �1t�|{�L���ܮ�������V~z�Bx:�B�O,��ӴW��_L�w��&<�����iKF^���3�q)gPtxpX	�W�����]��t3q$�%��"���E��d�by��ؐ��XMlpdLd�����M�w������`݉�pk���O0$:ε�lO*$�52*K;�da�	5���W9@�8.T��L���,�Ԙxݽ��J��s���9�q`c ��|)d�uyJ�aq��}(,��Z�B�.[���k���ap:�S�� Q�	�x@<g��j��B�k��q�F�v��9‾�ס��W����ơ��֔>��ɚ���W�m+��i�{�X R+�dϞN�a��u�i���"�m7��8EGj�;�=}���c��ֱ�eT�=��������1pJ3��k���/�#�y[j�1��}���6sh��E/(��z7#�!DS���,	;۾Eo'������S��Z(��bOFՕ�b)z%�OΖ�lD_�ʤ�íA��遻�s�E.*:�Lr,��������Ӏ��1K�%���I	i�H0pS����w�1�^�jz���cNI�}_�6՛4�ڮ�{��:��Fs��r�v�UB)��8	3���*����y�5Sa6�f�zdC���#X��<&���(�U'��O�X�۶��wL��l|�����喝}J����J���] $S=n��#��⸸�O�ՏC�18u�4�Wk�N��e���V'���ʜ��Rԋ�6�s�n�}��Z̀x�b�<U�<�a^i6�Ro\َ�Q�W��F��ң�m��{1h�z��,�譕���y�:�W�
f͇9�3q5���7?4�)Wrzn�9���2�9܌a ��!�`��N�kܪ@Z_��4a'��Tnɦ��8�rr7��rk@����{���S��Q�t���d��b-,|عVk�gH���V��(�E� E� �dG�Y#���e��Phxaz0Nd	ܐ�B��W�j7s���!��m┧�;�Y<X�ZI���(I�9>�%�+�"����$C�<�Z��l7F\c��s4P���H�.�v�R�:1�)��g��ܸ���7���5�t���B���a	I��>=�LH�kȒ���mO ������Wf͋<����7��RS}s�>PK���f�f�������J5Lx�oU܁�-d�!������f��Uؑ_�Ĥj��P�@�ӳ�	�����w;;$ ��Zc���;0C���#���&QזƲ,�i���6�s�ɽ�0��l� �8xA���!���J��!�R
z���IVkf�Bxdp����Z��*m�Mn�q��m3I��E܄d��9g����P)-�&��o�F���v< �����-ڜ�j,K�o��f�����ӟ��R�Ʉ�v��/�H��P��]vEa���w@�1���d���N��Aݵ���*��7�2[_-������Q��� >���\�a/ e�j���f昕�̪��j]�v��@���"���ù���f��Z*Ǹ���I�/`�,h*��w����'�?{��l(M�����|�m��5��j>9*�~( (���洐8��ƨڥ����rK�����h�L��;t�+$��s�&6��=ߘ�<�ig���P2q̩�
EgR�{�ك���+a�����"�I�"�+�#���j<;{T�Ժog�Q�g&�;�=�xp���L���n��L��M�I�t�y�����4+��y�%�1������U�Q���Bbr}�O�Z��g����'��R 84���b!qG+��G{�AP=�cT�� Juۙ�Y"�n��@<hT�Z�PF+�'ڻ{��2g����鋿�|���V�e���0��x�̥зO��T��ل9�}%�4�����V5�D���e*�� ��%���c��C�(F���9��R[(��0�
E%��	�[��(��H܁Q��ȍp��r��HYyu!�ϽGo�w�и*.jfv�`.��Mw�Rz�J96������VH{吀9;p��]U�J�$�s�������'�`Xrq��j����Ocuh+��Ɖ�/Ř6��F20}y썇&ҭQ{y1�V���.���[L{�����.v' 5��4�R����vGj���TiW��S��1X����=䚼t5�D�s<L{]t���6�Uz�Ա@�+�A�.3�z���2d���` 7O����wT�-uH�m�oQ&P�;T=㫔	J6��AA�(������TZ�-�d���w���<{:��G��J���D�� �{H��"iw�Y;]S;Zw�L#ߤF^���J/8wΎ8
����;PҀ�������t�/0)�OH�U�a�ƛ3��w���'�P���y#j{�@�"A�[Rv�6y�x�pi���͛{�{�O=����ARh� q�"���߆zzP�~*��7���L�.�Q�ɻy��@B{x��{e;�6� 	�+ȇ�����1y�ǣU��KT��������UF����-����Ӎ�"��ԚjV7��"��^�Pm�]���-ֺGx>���䮻)R�k�5@b0r#'�!څ����V+��YO��Oր��t;���<.�¦_�_s(�^b���H?����L̗���T�WA:�O�X���^�A���"�Kq=����W�o��sf���)J$��>ٺO�t}Ca���Q�W �T�:^�e��C��jRq �+j��f����7���^ ]o��^-\�\���Y$#f^7����3�~�&��y߹R�J�C)>�n�ut�0�:�|&���[�Z�y�!����ݤ��zώ$z�uL��hH�I��M<[-c�`${l����-�Tz40͟;����x���A[�U�S=�l��P��ɷO�@���tqCa��0l=Kg ����Tj.S�l��2�[8ܟ��L���v��;����!���Z,d(�wp�0Η|7P-l��+�d��:T��̲�9RB@�)O�<9����i<î�s�je�l����?��h����,TK��H&��n��;W�8c��E�Gw�uI���o)Tg�#F�N��L �l�2�gN@I����k��շh�U�B��1�}bN2W��!�(2S���h�%�o���;��3u� 7��� %'z<�7���#Ջ���Qb
�z�M#r��Wʫ�(������e�A�klׅ�����E��S	]7����ڥ����6���?!��g_fҙ-��ɇZ�imQ>��ZE�h���ZŚ�\j�͐?y���,�
�)�{�����p�Yt����L��SݕO��z��t��+��K�N�+�y�����]��T����݁"�vsm�S�~ny�!��&��v�\`��nyV׶���)��T��&���w a�C`SN�݁� ����D%{���r�D
�B:Gꮁ��#tsG'��@?nL�wS��DW7�����=I	�`�'|���|��bAa�'Dm1R��$ٷYl�{[��?Qa9E����z�,Ux
��J���$4��ѢPy�������Ev^u.Ε`o�= �٢�or9ݰ*l���14���F"̀K�� *���>�J��L8 ���ѭ����3��u�����Zk  f�+~������[����7��ס��|5��z�8�JW�a��;��.�H��?��ַ���W	Gѽ~tcC���^ο{w�*b��B�LB��Z�;�"Z"v�}�ߕ?���Z)���2v`��uw��h�<#x;?�_sY��"�Ě{�2h<+9g�I[3�w���A��n@�U#Q�����,	6"��g��홱�a���C�L75rX�D5�y�dV6�YCk0T~ �(��5ʡ�I,�K�#�X���z�GY��ޏ�@^̖B�z�g�/����z�=l�;�Q�; I]�J��J�[��q|��G#����r�Y�L�Yz��5�?Bo���V8��լ.�s5��_�1�5���_.	�����r����Rbx�vtAf	��O�˨j|�GD�!�:�s&I �H�x~�u^�����3s�\\�ʩ������6�� b��U�Q]�;>�w�Pe{��kF���LB����'4`��(߈��^�N��.��շuJ��J����r@�!��"�{�bЈ ��"W���C�!C�������$�)�j���酂Ag�H�c7�%P(L-.��.D�����[�O�u� Ѐ����֔��� �Z'�͈�`�$�1P2z��)8��r!٫���������m�.���|��$�� ehJ�Jg�?٠��3\y��q~Dz�`6��|�\�����Ly���M��v�(�q�[��t��O�1��7Nf[����:'�vb0
_���MՖ��}%��d#�|�n��hC��oFke�XiFk �s6/.��x�:-Ƭr�����R����wl0��	%ы��A�b�fJ��@�Ղ����u[�Q�^�p�Q\ͧl@�sr�	A�&�����=)%h�}vC���L���}^�y,,K>�[2�?��m%�3�y�,y�@.������c�~o9,��x�紀����(	Řa!�I�?M(
ܸ�rͧ�;��Jo$9���d{��@ |���� �{L!V�Q}���cwv�<��ӷ@��8!T���T�j����t�M��K;�4B�̣��"�HXn��I�T�q�������bzoV�?�O7�[�%�/�,wF��6��T�S$�~l;B�&\Zi�i ����`R�u�-���}��̨��u}��&5����� s�׃�q%���DG��W�y���_1OC�)jEK|1�e)����C�֨�sM5�N�ϚZ9�[N���A&���[V�^�ؾ��>�f��(�e����$y>��!��>p���2���B-y>#��R�⟽�{MƋW�p��957"����T(1˼�	m�:)H���$�R�.�v܇!��d�PP"��'$ψy��R�r�n�v-��|J�	����)f������eAxM��!���ԑ�v,'\�����p�IQj>��$���L%�;���j��W����x����`��݇*	�L=�{����jS���ul�ѽ4ԍ�8�ʹ���5бG�5p[�c�n���(�24�ZL�515��_C��\�O���>�7�)�KqE��9B�!���C�#ztR�~�T�M�63�8�;E��t�Sq9��A���]�tJ��P��d�ߠ�~�����
��k�T��'��B�_׎I9<#��z&�Zzb�9m��6��`���R��w�2��U
�̱Z�:z��&#����V��u�
�9����f�<֮:i̜MV#->n���<*�
B�D�<��c��E��w�C�[rH��:��ٿ��(�.܈�87�.)x<J=~ǱZ�V.�oK�Y"Ǫ�_oJ�-�U��Yw��"�A��!�+�r�_�"�D���1< �H���&���7��M��#�ng���ǉ疴��@2ZV�_>����-��i��T�`㤯�g@�{��S�s:!N��2�V��@���؇�F����T>��'5��ә{��x�(�p�i�D�.���f�uA"B���())L�a���+U��ے�#;z�Ѧ�N����:�!mt�`��Q�Y!y�I�bpJa��I���z�a��"��<q�P�U��d ����hx�S�S���j|p`%6WP|�ƕf<O���ܙ���k��@V8ऩ�G|/���ϔ=I`�����3Y�jÇ���A�9��y=�E��	E� ~\�F�>tG*X�մ�~s<-�,2^��A���%��C�d��*��Ĝ�ڟ��I��z�a�h>�@G]��NA��F�먤���%���U�04��mC4��CRS�|6ìL��S�Q�.�QpH:y̔�?�d�7��5x%��g4�k���\�� $�E[X�|�4$���q���Y����e<��|�u�!8Ź�%Z�+���g_�������rS���\}C�O�3D��� �*���?����y���/3:j�6��×���M�,��>�,����E�T_�p�7���1�Y���&B����Ļ�)�ޏ�Y���JFz�_²�tNǿ	c e8�މ�f���!���}�y�gl�����1�Q���H�I������5��á�i�F��ijr��L����)�g��~��?<�qD�(n"kgx�w�BDx3V���/행��w�E����;Mk�ø�kx'k'ǡ6�@#CtFZ�e�>���.�w2�O�=O�턙�6�~'B�)�u���=f�Jg
Ġ��r�?9�Nf�[�9|��G���k�	dt�]�܄��l�B�oN9�VL�_qs��w�� �>�v�k�N�R
����ϛ0��O�m�ܤTٿW����~G.M��F~H_<�.�9�$��_�8V2X'��l��8�;�Vׂ��U�M�Z$��� BR��N|�Ì��ү�О������~Z=G1x�+��$�Vl��a���5%���[>M����ګ��Ϭ�;R��+DD��� 6:(W/�e����,q��� ��F��*�g�����A�wS����C���- Y�x4��-�	8��o�9�d��~�)S#�7*��0PAX����$5��b���3;��$����q��l����!�@���AO�P�YLg�˪��,�l�$��<h�Z����邌rP1�Ա��g��	T'�!{5n��=&��Q���@i�XϳRV���+8B�Lڻ�a�3j��ҧܓ�*����rHꏯ�Ƴ����%�YA�mǗ)Kl}ξ��V:����m��ADR�pN��i<���&~���jn�,��5}V��۝�$5�RP7.�d*D*�&Z�Y�V/Om�V����� ��ҧ���]��7$�}��hQdN=�Ɍ4_�B�>�g���ȑ9�t_��	�wC�a]��~$?��/Jl��g�I$�|�kU$�k�`;9�̹?z�l��ĕ=�`�Mt��E��G�,���+�C���-B�{�)�c'Nv�O��	Q�=f�~%�,�c�o���vb��+%��	1�_aّ������G8]��Z�%�O�:�S�@�u�ͻ/�*��ʏ�N��7�i��������?��X��д��|U����!�5�71^.41[F!|�ʶ��ݨ�ٔ�7]oJ_��r#��h�3��Z�s�|����#MV.��)N'���Фǿ�]��ȱNQ;�{���\�����@�����,�>
¸�S��a.�ٳ��8��/v�t�%�Uq���a[��1�A��7��r��¼!"!Z�jUV� ��@�դ*���"c|E`�gR�WppX3�m?e��s��}Xk"?(�Iq�O=)=�h[̆�5�pM�f���Hl8�Q8���;Z�1o�v[`N�O���00pU�F��Ǘn<��D[?SR׿�a=b���I�C�\Ɇ��'���B��-P�gʂ�1J|L7o{i)Pۖ�2�
��8���DD���P%�Տ�PK�o>u�y̗uL�-Ɖ���W9g��S�_Јe�o��s� .F�X�v������b�ǂ���/u�����ǽаS�d���X�8�wؘB�n���)Jm��éP �qD�DC�+"C�vt������}4��	��AV]��H��F81�7F�kB�x�x�Y�鈢/r�:B[]-�[�_�3�v:�-`Hq�WUۣ"�:�s�=�d�������*�;��
1[���[�إ ]Մ�f9��(��
�vE\Y�f,i@3ۇ�==��E�?�ߛ�Es���jb���F�q�=0�҂v��r�ľJ�B��.��8�E��.
��3�5VUp�h��vtA�(�Z����}��//�|b)��ij�P};�����feF
z����w��Q㶟�Uu�K"1�=h�5�޷G���}r��G�߰�^�t�|r����If��č�r$5>K
z�B�83�r�te�$�ב�5�N.m7����11�H���� ~c�j�'�S�-�/F�wP�/M칋���nF��Ҵ��GmB��o�kf����d��������(%3�7%bl6���42G3&�,�@'��C#��Ң!��m�����/�c��Z=�����*m�,�����Ü�T�[�՟�,�sϓF&_4?"�z��+�b�¡Yfh���6�ڠ�U�zO4�yt��#d=�A�H�"jvCNJ}��U{���PY@�n��+v�^��纴��	8�3�]C�-s>��9�,Ɉ�E����3u��>O�WX����{��r&q�pݤD��p\��Zz�?�E��N26�� �!���gK;�e�!X�����[ �ap��(��9��Ei�8���a�i��T�b�K_��"�y$��l���ڑ�E���>x���.��v��VUIW�b[L����{b~|^�i~%�5���E�Ca&?L�b60� -��(���+��o5��N�㇈M�b�ql�|��-��f����/�)�j(�0�h�
KOH.k��o<�Y�4���c�2�E�Ӊ)�+;�`�W�Ѵ���س$M��Q���{�#����U���[�EH��X�#SO�5�+�dh����5M�U ���o��s;Z��_p�[C=@5HԢ�<B�ȵH��o`"Yx��:�����>Kv�Q�?�ʚōG��_�)��X��\\ZCV�H�����Jf9�$GI�P�X�t�<����Eƻc	DF�FC���"c<r�{��~p1�-GTbϏ�ճ��
���G' � ���]�(���<�"��/�0��^N���/��g�M3n��bD���7S��z��pNߠ�$1q�}��婧����/��=Z.	��zl�.HO��S8
�l�Nf��:�
oWj �.��P�TP���@�r���LO�88�t
�3 
�g���cbH�	�����|͡F[�^����20��S�&���=
Ʈ�튣.�ip/O�ḳ[d��p�j�!l<��EL3��@�����p�i���sګ�ћ����+���j�J9��<����K����?C���$0!8�1B�����b>��C�(�������O˙HP�v b�F�W?��2��L�Y|Ra�)�.`��W�����:k�J��k��@Ƥ�z5Ҁ롞d_�� ��r��#����^O���������!�����r&�#j~���-��^{R&���ͩa�3���R@���n`��F��DAJ�lE|'b�h��]%�g�ł�w+��!Uq�>��>"1aVdb�g�i,S����~}���I�f�X f��1��u��J3Cr.�)
�dT	:l67�h	�+�$U�x9$�����3�_`Ǆ��x,=�]̅+,,:I���,�_��oN�ʃr9�<��-���� %���%N�I`�D�}/ Y���ݽX��d����"g��vp48R�w����h��Xk���ȪZeA��p��U�
�Eb�sC6�J��T>�5���7��H��7�'_���?�T�̠k�vT��!�mW�o_uQ��2N��v��=]d��@|K	\o���@~���)3I ȓ6z��Y���"9h�ԧ�n�9�܎=ӫ��HQ>��_���WJ?�ٖ�y��\��U��Ӹ����.�Nh�JjR���]r�O���$h�=l��|��g"����V$[��f�,=���V*�:�9�����]��܏����%��f��~�վ-��v��Ŷ��hĢ�uN�h��ԯ�d5���* ـ�7>x_��������o�79�9d���O�W�6^1߄��^�"���=2��Y��=�䴧e��M����F��E��v�P�hj,A3����̽����>����RS��2�c#���=$�a���ۋ	>Q�e;�kڷ��9P(KW�����KF�apP5/�3��F��;��y��'�N[��C��E�U����КhpSg��z+pٯg�i	h-#�֑-�H儸%R��e�ff�5\>��hpn{�[i�ٰ�͵6>۴J��zn><E{�U�?	�$�5i���-�#�lC�ιݹ��b����	/���V�J^�N'r��2]/�Efpf[�V���İ�=��W���b��&��R?D��o~6�<2(��Rkm0�ȇ��@5TLI�v�@j<"�s�L~]�&� �ȁ�+�=��ʃ��31��侽��6��2+�$�0Ĥj��|�r_�9��sO^��m�ˉ����ϽD�@�՟�0���ٓ��:��G�SlQİ�Z]m�9�x�"���/wo��{)�@�1��\�B�����ٮ;���fw\����vu��E`�"e~A��7Iu)�<S�'п�x�yJ���� �'A�]k4(c�;kG�b��N���i�
r�񼹂�XE)�~���\j��О�Cmq��f��(����X鰋SΈ�B�E�O ���� R�qF�i�#8DdȞY�xj��	Di��,�ݯ�<AƟ�5NL� E���n����I�Ժj]в�f��.��R��0����H�)��x��Q�d�>�}gͤZjs6b J�g�/���h?���%͘7��}�EU\�� /]���c�\�;'��_��;�3�i�D�|��]<jii��A� �]��d��xY���n˞���,��kj2�Z��yiPs�7�F.H��Y� �xg{6GF�[  +��`�@����ʜe('����L�CS���㮴S �ao���F�Gz�C*��X���l����=�5<E���xV��u#Ok���>�@��S'�5�����5]�� ,|�5ߖG9�-q������y%��1;<��H8'��}�:��b�Ư���8h�\��8�ހ>�u6�|��j�:�}���2U�����"B��$NvQ߄��=뭕o���̤
�+i�Tw�9�Ω�iʚ��?��'g6Ղ�������ai)9����p����o�o�V���`��&1ù_��N���w��d��Cv��x���$kgrs^m�m��-��XhҬ����^9�i�I�8xB���`����4���&�:cw���G{�Jj4����.$�����+*�A�g/R��N$j
[�kp��B���n��j}�L��&�q�(�59�\^����|�eVN�hׅ�ǐ����Eh ��$�(T�['[�~7��"��,ǉ,�p�ݢ�?�Dl�|&"�9�Մ�6Ha���Q�ﱹGG�s�#������g�$A��ya�{]�߀�uk^S��*�?%љށ6vr�=LQ^�	w�S{*�>i%�G�s��#�O7R�孌�x�h��f��$�Pd���I��]`�P��s�*V8@��(�����!K��!�#��r�Aç*<�Iu�+�<9�
bQ]y�W5�������N�)�rkM]V�L*����.�	����[ƞy`&P��Ty$@E����:o'H� .4X�ݓ�KH��0ڄR��'�n�'��Ӷ#�L���$as���5;,�^��s�M3��m&(\o��3]-�`�6 ����'���4���ˮA���`TU�M�ANtwU�p#�����4m3]k�E, ��}�=��4���0L��q\!#����#�U�� ���:]�u{���t�������V��BZIN0�^��U�Pc�(=��8ظJjg�¢�uA��2+�t���W �k}�7���SAVtt"7�m؟�C�ǵ94���ܚ�O���[��R�w9N�ht���
߳��Ò��Tt��TҨ����);��?Њ.���.n���0r�+�g�>'��<Z/�O�g��&")�񿒺���*�Ǝp4�K��>za�
Q�=�|�/Xz�+�DZu�XKX�Ý}j��/�d7��$~��֍��Y�AY�0�*VP���ȧb`kP�W^���w�Wq�wE��B��MlM��s 0�ߟTH�y<tV�Ы8�v/.��5��9i�U�I��`�pou�\�!����g�o��<m�'��-�[���ݕ(Y���'��Pc~b������f��_�=�D���+��Jj|u���jٲ����h1�CA� ���7F=Vg��S'����K��﮷�3�O��z��aN�L�3�6��`N
��r�<���n7u������.�LQ	9���o	�^�����K�!H6���6�!�ǘo'>,�}��6�h
�ݶ�熜t���=%���݃	-�� IB��9䀡��b�zM�K%��'��Maσ�����&�3�Oe��$CN7%��}�[�)�] L��&N�����
���� n[R�3���"�S֧��T����a��p*��?Ik|"Q�@�w�ba�����b�~���[�G��n���"��0H.�#�z0��w3&��U�,9�Q��.U��w=�\�]|�,��5���3�,�h[[f���w�9�k�Ǜ�W�@-y���823�b{��S��$s���*�:k���U3j�cG:�q��+Q��۽�ݲ�\L�����D1m�y��"&]��Nw4���"[�>R�(�|�ֿĬ�<�M�
��u	*�n
�7�u'�������HUjUG��6E/�wQ��a��eK��E��3Z��sk��P=)@�d����xf��U���S]̴WE1���Z� /&O��Ht���xz�,�l8�J77=Y�����u��7n�Z˥���d�h[@�%�m��h�O�}o=�U���˶��`�J���~d\�����o��p5������aC`]5+��B�7j|j~��&|4+<��4�캈��n�h��GЦ�l�2��ɟ{Dg�aT.d���؁b?K��9���9�G;��q"�l]H'>�GR�q+��5�vy'+�
#�n�6Mso)j�:���8���D�i���$�ڃ_c�#2��*'���ҩ� �S'� -�03��q�(��[�`�-y�Js�-�,V3�
�wh�}�a4$4�V��;���ѻ\�j��������)��
I��Yw+�$�E8���Z+&0<?���Ǔ��/9-ӈ�9����xצ��<�pC�e�.d�� +�ˠU3��n�w2�q�c.�\�*���`#��DM�6�HW�c�8���M�"=����հ��T��i5�������3Ϊ)��ym�M.du�T�KG~#t�?J�GZ�7:��$O�0�f�C�������}E��DT��R�Q4�Ό�p'�)C)��l������7זk���f�w�I�"�0*f2�o
����D��G�`+__V��W~?)I'N�J�b]j�Lм{�A8��E�]]!�'+;�����ה4o�TRvcF*?��Y>E�5�3��֙�����d'����ǖ��Dx@�c���i����v[���>X��D�`��j�8Y^��4`W�`B����ȵ\�/0��D�s7to�i?)N.��n\=-Q�.�4���`�� �nń�֩X��K(˷���;�xI��,�ٿY"�������Z�R�����|zE(4]o�U�y���	���,0�Y��������tȯ�cԚ���._�~��4w�#X�q��|ș�Osv���L�B��j��w�XQ��~�D�'W��ΦW���!�J�3N߮�Ad+g�у指3us��ڠ�	�a�K�"N��G�IѾ��j��vԔ�5%����h�1�~�#�y�B~<���Eye�{{K<��=�Y�Y�8�7��b��� 1��Sf�N�h3��8��dgj��1PQ�����(�cE�%�`�cwh4�d�R'x�b��ǵ�н�g����;��a��L����H�]Gm�B���pg4�>sƃ����y�Z+���3F�v�P�D��ժ³�M�/,M�n�$d����]���q��/��0Cz�g��xcO|��Q�냔Bz�uf"+R3|!����UnÕ�u$���3�(N��h��ŷ�s��p�B��" 	�Vj����1$�#�{�jn'�f�M�$��"���>a|W{�����ô�i��1L�-��J��<
�a�8�E����_��Đ����
3��K(u1S?�N��5(W��d�}�_�E����>�|?q @�m�sFY����}m�����N�9��ٝ�oO�'��,%	T�?�+%���<���܂ ��H����X���'�}���L=��9�t�g�� +9�*H<F�rFS���܎L�?��Jo�*�y�Ԡ��f2�̢�_��]����(8��s�*�8�FH𭖡�gB�!ɑ����N#J�
�M������X*�ŷ�
��{�Y��VvȐ����4��m8�%S�t*=�~��[)i����D��A��h�0w��娞ו)���E��HL�5����Vk
� .��;�W��u��S-�;8@e6�y#�>; Oh�u��eAV�d(|�����2�s���O�C�\�J(	�1�v��b��DMy~A���,���³�?Y��s�z�i��҆�K����\�N(���h���ۉ6�A�eL-TCP̣�	�T��+h��c�� C�ˋ³��d���Q��j�ݞqt�nP7��Rm<+:�Ol����,�b�>����oj�e��˽.#'�G�n	�8ǵ�f��Ok�k���!��A��fPD����o�fLc����#���^��N�?��oNv����G�G#��:U�OHw^�����>
'��W����P�QE��5����>lw;�'RbQ��=� Ӛk(�)�����\%�Si��JH�'�����tk,[����wє3�&�)��`�t�B�k�r~{��R�"�(+��q���HA���ۥ�M���C��)�9A�2�9ErY����
��X�@���\h�D�-��>wb�uO>t���ǳTvQu;%9���^���@�� M� �o
eO�RJ)~<ܗr5u�q�MC,	�M�PK'�<��	çP�$�-�kE���YY��������"���N��#%��.�I3`�	�)�{��_�������i���8�:���F�5�8 @%V��N�"B�\OrT�J���uD�P�߯%�cȏՉB����0���7d ��@�k��`|'����:�)��S�����Vu8oc:�~Z��S�+Y�RC�
���^���������ӓ-.�3_Y�w9�	�����c
�b�nlZ@��,�$�:�	*�BA� 	'l9����n��`������C�	]��_e�4��de�
����5�c��J"t�՚z�1��/�bPه�A���v������c�&�A7)!���g�2������Bh��~�r
�� �������Z�s���=p� <���|�7��a�d_�Hc=Y"�qZJ}�S�By���VS
�+�֋�:�^W�ҟ�)1U�k8^�Qw�gme��Ԟ�A0�7UӦ=�+�C�6?���L�3�:�\�Aa�����NL/d�:�@kZE��D+�>�E��Kc��%I�B�z�շP ��ȕ!���*���q��_�F�{w7�z����	{d�k�|,�NDv���"�v��=q��WR�����NF��S�"�������Ce���m +ے���j�����?1�ƶ�����>~IE����ii�}^jqߌ�ph�қܝ��?�n��&�%�<3����uْP.��$'y�ۀ�	�Ҽ#�K�X�߄�#�ތ��넡w.��1�M}W�]R%:X22Y��K��}�q�ϙzw�Z�V� �b�b�D�졞��6���1��E)j�c a����<��ku0!�6��:7�hr������k �eᑿ�<&�r�TeW�k�ujb�PL���6'|�[��fށM��p�Ù��>P��	��r�'�,ل�	F��q��u�Fo���'�2zcGBtC�݄�C�γ�?'λ���H8�-�;�)0�Tm���_�\�6>���ȱm�:D�Vr�럯r����Dʶ`6����� ��n��J!A�u�!.�J�8��g�شg�<��m�o(k�Y�;��c� C�6gxdεI��Z)J��4��m N#"���;��m��%��9����ڂ�.mG,�0���Ma@i^�_���,�͡��b�0�n��%�HkGi;,g����7	~�xh���n�bU��g{i�n䫾o$�+��	�&âȢz��,n�8膌Ѓ�]JC�'�$�� �gW�n�Hڥ���V0Py�Z�q���;|�r�;�X�d�VPS��)k�Hu��Ȑg[�FcS�e�/Y��|)��l��J&�s /fZ�|/�	����?s_�)v����.�+��b"��WHP3�@�ѷ���p,�}5G5��g��˒?vha�zW<V�C��?�l~��������ȵ�h�Z��+��Lvn��8�O��Mvi�е�	쟃?�J���������CRN�/��$f&Nw�(��n�n��%�أ�z�.�C%̗�;R�ڕl��r��|@ ���11[��D����om�X��M�Z�(�p�S�E-�u�}j-���@�]�{E�R$��+<K��x��/��O�s��K�2��G��$�-�w�F��=��v.�����6�j���2���uT�J/t�V.,b���|e�I>E�]r)t��*��yO����H��,�j�uS�T�#��ͣ�9��jg5�� K���n��,�<� 5~�nR�,��'-(�R��y��Q� �r'Q9q�
%��a���P�V�@�����`�x�\}�����wW�/�\k�</SN�~ȵ-�p��#�2��1��TN<��a���J1�F�Q�=�g�e�,��
�@Xش2v���W����ڸ�~h���2�"NN���� ����~��뒦#�Ȭ�c�%�qq�?��ow@���L��$�^H��(�(��9�Iǫ��˾5'�� ���o�<V8x�m�5J���W/�ڦ��b�s��'S㨅|D�(�J�	�;�U����_����lȖ���k�O��?���)��Kez�����ބ?�\��k��!g�
����^Յ���Nq(z�b����i\�4�\��DL��4[�z�^?UQg�(����B"@���E��g�Ǣ�^������07,������|5��=��A��fu/�#����
�o�j2R6L�H��͉�gR���t뵪PD���ŁR�otř�On����ffz=Ԯ���ZNn�o�8�MB6e:&��X������xP�d����b�V�f� �ޠ���AR�E��w������5��$�c��ބ��J8�ԣ�j����R=��%O�f�Y���>�O�s����J�pa���T�G�ϓ`P,�Y ��ȒO,3����l��`an��m�i��)U�T���`�ۋ��/��*���$j����}5�Z��oP���M�-	J�B�SQ����7���v��N�R��)��QF��v8�v�c2[$����������w���]�5N�)�D+h-�-�-bDj'�
��٣l�xK^r��Vi�OKG�N�H/���%V�*U2�JX���L7�cU������� q��P�ƀ~�6R�r��;���'8���&��j.�����x̭�w>�%�#\����j#9��/?��n-@栌�v�����҄�+������oB����th��z�h��5^`��iX��H�39��g��rt�E�/c�n��Pn��Te%��K_�]gA8�wI��Du>�!�A�x���+˫��tF��z)+@�e�_e=������6��k��a��MM5��o*�1�5����Y�����#��hsn��,�xx&"8֮ �Ȏ��*�7k�����,�i<,���/�4���j�v �,����X'�+ю�Mo�n�,���>����Z���Cd9Y?��|Z���[.��	V�ٟ�,�S�[[je��?^�"�@gq^^���#됌o��)B�|[F�B��lH�?�9ѣ�F\n�?��+/*�c�^�.*0ퟢ��֩Ŷ������o:fh��U��_�M�G�G2��BA�@��r-|^���Y�LU*�����Ԙ~sWrF1��<�f�)_%
`=�᥂��ݸ�����dZ�(W�x,��ʌ�|�"@T��n�"`�n]ڱ5$���]��G�$�.��v@�(��i0��Ưq#IS�/������J��iVߵI� �Q����������<_��ד��ȟ���;�n����@W�y Y��J��X|ܿ	��gZ�Ь�v��U{�Hq�J�4_-��F\���޽�J!����]��x�D��~��d���L鹐J���Q$�Ј��3QC5�v�"VZ�r*G�hAzԜ�����I��,�ie@ݷoD��kי��M��RB�ĿGi�=����[�=XZ�ng�v��.�xﰪ_2�.����1���4p*�hzp����`S�me*�2�Y���]�~pj�Z+�J�H��,�M(]�,�7�/RC���k� J�=�5�H��8}V�P�oh�l��3����_D1�Mŀ�s��ϡ�ٵ�Q�/5M�n�
��GF�����b�8D����CyU_0�a�.��-��P�'��/l���Z7U�\��v��Aw�ՅG�U�� ���gs�uRi56�dI�M�JS������T*�SP��� &	?��:�R��3�Lt�\���>U�+��qͷ�QS.���Sڿ��Yh�J��Kmt�%�uS?�d&�'A�Q��)�J���er ̚x،�@�v��gF{~ ��x��ͮ��!ir�V���V:]�7�G��F�y%��GZk5B���j?:��oTR�
Q��� n��Q�X4�_)�N�7�O��I�0Y�Kk+	��J��>z���[T;%u��
�x�ؼ�U����d0�pLum��	���c�g��Μ%��Y��0+	�RV#���59����'t��,�����F	h�tE��D 
��f*q�![�?�〮g������b�h��^�x=,�B�C��隐��n ��z���g��Æ����q�ħ<@�t0�rԑ�Ӧ��v�c����v�o��U�����UϽ�`�C�D�~#޽
�{r)}dn�"� ��j�Im�Y�L�%�Ҫ��/�[wN���u$q]7���J���|��yU~���
p�tq��&{�3Z����\zL]٨����D�S��`����o�-ה_�ڦ��+B�fs��"�Xo����mԯT+>���KЈ;Y9�Lpb���!	��)?��{Q�#����ٱ��c�â��/���?�����̠�������e��->�^�+���S����]���S0L&�f������v`K<-��ڞ�;�S�#cG*�JQ�'PO�ZR�\�C�M�E�v�G���įz�ު�{/��$��`���N�k�]������$�Gb]ɕY�.�@\���.�PRX�.ؽDԆ��WK�	���zm�v����J� ��!��2�+���(���rn-�¬A�!�J^r卑���j��*ԏ���,jɶ6���58[�R�v�z�i���p�1ڸ߭'/�H��1Z���K&����V� ��.���C��7U��'i�$,��Ra��XEr^��!{���tLě@�=�/4�u��Х��hE�m¥����o�yW��Y���3~��bf�g��O�T���5�i���K#,�Z�X1z��� �G�����~6ٟX��y�b��Ⱦ�>^�\C���hrN��̒)(G�]��x�ܴ�����b�!2M�|�������-̐~4^�@m���ц�����|��f���W���p{�z��G�ywN��H�ӧ]^w�Ρ�O�"�*Q�R�};Kv��*���'Al����Ț[��� �=(��tv��"�Zؚ�5T^�������u �4=�F�B�r����F�	�u����3og�����$���c�8�"��k}�E���b�%��L��-&u�
�/
� ���Hq2('y�h\�1�,��(LX5��ԁ��K�e����`�� ��H{d�c\Ď�U���qg2�]��`�}��.J,��R�=�\|�#H��i A1v�?���+�_I��m��˒�� ٍ�lHY�I5�Gzƺ�/�a�!����tE
ˌv���e.��Ğ���.n�*jO��5�6�^+|{�$���L}�'&�ЂC��m����J ,�L��/���ٕH7B�\ h�P����
e/7�G���V-oԂ>���L�L�&��b�}@��Y�&��J�hsm��o�;�xMt�J�ұ̷�_��QxJiY .ӆ�!�YCi�B��y�.��|�oޮ������(#--�^p�)�u_�mv�ۯ\�S���n����wo�6�	l��X�D�x�$B)�g�qdw�p���#������'e[;y*'����zǗ}�t�QSe�#�&��kl ��
�Yeh!x:�L����mNPo>̭�J�fhrA9ӣ���d�!�h%�-.� Ő���'��}�Ѫ�Z���^��,��fr�������� �ZH�m5] �a�cjįR��k �WF��8ܦ�9�ݐ<�C?_���VL��_i�N^H���c�GN?��Q/�qZ9���D�^[�D��8�#����h�"y�}nH��k�C1��z�yû��Y�sR����nІ[��&6[I�w���0P��h���/�=.u��=��̳C@�M��,��0�(B1X�����{JLX���H����ܢ��v<�N�u��&�S��FȮ7z�@$�v��t��aҖ��6E�1�P�{(�C�g� ��gg�F��${�p��M\(�tjǹ���tW9!g�Y�H�`Ҥ9�����*0�xY���t����R�k$���h����F�3Zl<��Oi�8j�,h��{y�h��7�{�pWm�Y0���BN")��,�"���)���Q�H5�Z�l�;��Y%{�qL��K��Ҳ�������gOKʹ�Z 	_L���F3��y��J���]s$̭.������� M�Azû�i�	@�辜w�ĮMd�X��11��?��;Q��IG�T�O�b��ک��ʫ�h����J}�>��\��� ������)  ��Rώ�2�MS���1��u)�j��qá�¦��(�GK�Z#<��L�륳�4��<�(�N[_��|^CY�ok[��O���_R�J#�+����c�EK��������V�,�;WlQx0(	�{��
/��A�hF)NhS��	Ά385��� ��l'�τ��hU���NDbĎHe2�X�X8<3q5��������蒖=~�3�}
�mv����|����0��6Dl�1W�f8���a?P�3R�**��4��<�!r����1�Ehi�R.�T-�p -v�~�O�l���6)���H��l�����%��d���\'/��ݲ��U�>�@��!�ԏ���w ���GD�Nǫ�%йe�y���M����M�����]�~�h#�$��.�(�[��Fm��'Z�\ԺFMC��_`��jwF��m ��_"=ϤY; !G���G{�NY�w9Z��XG����i��m]YB��#�\��]��u��u�%w��͂1{S�^5�W6�R
�W��Pe���m���PW7�v`__��χj��V)9�0��RE�� /�,�&��
��y잧���Y�VOb�ۏ��i�8�Ii��ø�����.y��M���M���<!{l?��J��#fT&i�3��WP}� A+A����]�=�oK~%�1(շx��%�+�������+�hV� ns4�[�' ø^�'L�y6��{�қt���e'<%��4�ux��8j3"�g�1]L~�`M�+Q������w���]Q++h���fJ<&�NI�d�}�����󛑛^ؑ�tyb�h��P��_$V�?���Y0�R��VXa�Q�P1�c���bxlC�
�P�ER���A�|hB�,sȸ� �����14|�[^0/4�j_���ẼC��eI��և��x���F�؍!�K���S¸���4rW\ӂVqyY�-���B����*>�
k�5�w��vX���'i�l`��+�p�!��#�8�	��4%���t�G!��o�x���)<VʌJ�M9�]�	;�;{ ��gME��r���ݸ\�NY��Ф	�z�*�l>�~�|�'��S�3�+��_�:ϔ��bvsݏ�ě���=bI�Nu���2�e:b�o��;� ��M�'���7~-����E���7��U���/�����wM���U�|�~3�����@ڒ�������*��/����&
dF�����3{(�5ko3����,W���&C`�J���)g}�X~`]h"�/A)�\	�E�k�	H��ZM��p����(��u���o�$l��'��o��o��i�)�d�?�GW�?cܸ�ޘ $ØO�ѿ�,n��Ĺ�>�f�N����"O=��A�z�o���r�u���I,cm�ZS>�ַ� �q$v�S�S�-W��T�'`D��wQ��a�J��|�IT�����XΈ"�{�>ZGx?���L��E�i���<� '!�`�Q)�8�iU1��9�f)D�Z�;̹�(�Q7�,��2O��ө�<��ʛRYd��w�p-(	BW�ۣ�~J%Y:2����/����p�)8�v�����.�fr-��2X��(�'g_(a&)��q%^
�5mG�1g5�Jϗ�v���ʲ�S0�m�I�O�PT�?�[�8�����Lx_���a��|EL^
�r�$��N?_��|���o��|U��ĕ�g� ���v}O�����m=�iTa �B9$C��9^q��ֳ^Q�Z���X7Q��lE
�ɽY�e�L����ъ��0@:+{$�����{C$����o	�;�B��F.�E��\��Z{0� o��|BS�EI������VP�E��5d�^�}�z=A�B�+h�.:�;HT���F�$�N�=��5=�>���2[~W1����Bs��bgƶ�i
e �Q�4�w1T0K^s��ޱ���m���?:�i�4h�-�2\Ƨ�w�#R���3lM�Q��tPeS|$��+�����#�^#�H 6}���L�۪1�t�̳��ӥl^�!���t���Ǳ�<y��K�`��8Aq���i�pe���xI\T1���G�,���e �]z�4yġOR?}��1����-���F��f�U���}2���_x�������#K?d�F�ౕo,�Fe�k�^˵J�fš�r��xH�Wh���_?��m~��L��X?7�L1��sٝ�P:8}��)���a�ɴ��ӧ��)M�nߣr�F��L�nw���U��-��ٴ���K3og��K�� ǈV�M��|�V{̱ɾ�])���Q�H�o/8�:��|���6u�U6����.��o�ڙ�'��Rq�W�I:ͤ�=L9�b[��&fKN����h$�1q��� <��a��Ӷ���x���6���~���j���-J3���)�x�,�|�u6�#aêܖMQ�i���.��l/�%���3�����Xۣ*]�y���L�����8i~\GK��;/��8�7����LM�Ѻ��[�<�#��3��[n�󢔖?)��."��D�c��-��*����@[�$y�pp>:)����h���j��1��P�����p��k��/@�����/����_Ɔ�>��d֚�'�}j��\��K@�7k��Q��{�����y>°Y{bq[�����r�^S'�OF�xY�]7q�آ����*��3M����~�(�M�`p��vj#)�u|�r/���A������j�c�"�{\A�l�����;-y���IщP��F��S�2�/i5����Ǿ<j`����f�rh�y���~0�Z0�K���*ݟ<�h4%5�JҽL�ʬ����M6Q�Д���}�Qm�=E�Tif`�q�
���dǾ�l��n޺Y�0N4KW)�yՈ�.17�oK�B��3~�UY�.�B�i��;���ʀ�!=};�i�(�M���w���\�kC#k�gzjr�Y��f���?��Z�ѽS`�e�d���F�����ӥ���ً%��]��@YB)���R�T���R!jqH��O�k0_�L��� �[L�}��)l7���+`�=�9���T�}�ԐQ[��;0��\H?1�����n$�!��<ퟠ�yQ~��	�v��au:�r�xʧ�g�{HH�F���C�,�� �m���+�χ�z��|��ȟ+$п}p9A�c"�+".�>�]:����';|.K8fvǢ}�� �͙b�R*�?A�kfJ���o��4F��a�������7�L�i�1E�R�e�� 6-��`���1��[�~���E���=F�ԛ������sm�xQqȪ�Gn���&�/oUOY!7sZ!���V3~Bb��u˵s1��S��텿�<�^�=�Q{ 	#�53�`��� ���Bè�I�x�O�~hng���N4z��N;��9Jt�Y���9��iH�-��-c|�I�R�Q� QN��*Z��u����VGh��� �����v`+����je\"�(A��5}<�%��ܾv6ز�dt6RטѮ� u�ш��z�~�W���y��u���RpkҽP�X�|kd��8,���9�\����/�}h�my�]���^�後S�/!͹p� ���H�F�F�y��,�3�XdVf�]~L��gc�@���������HP�v�%���c������ʐ�]��n�R�(s>}����^�q%Q`4a���o*Y`W|�ñ�=�]��, 8|q��Lu	��}��� �����u�\!Q�H��e���� �,�3(<b�#��K3��`T�bb��7��GC*j>�,�yه�IgQl�D~��C󷶧9�+��t�a��ܿ�e�D&���8Eu򀗍�,2��*ݕU�	=0�[y���wn�i��hWh|�W�ݞR?�]V�K�Y���O'�M$��7�{ೳi��8P������(�G�E�,<G#�/�\��W�'�-n?W=n���֚�i��b���X�G`2�(��I~��n늃i��E8#*�nR��/�v�\���)��8�����f�����}��1n �;wcDk"}���nWӺ8�T�.� 0�bT;����Zg`'��T��2�픗�#�4�S����ʞh����QK���):Uk��� ]yx����������6�7B���B��J#����i>78�����Q�aiȩ� l�� }��
 ���$����Pw�ao%��=�1��]	j̥��![,:7&p�r�(:��F�_ȏ� ��xX���//	�^��^�ж%|%����4��u��R�qS��y۲��A��\hu��8����e�IvVDQ��7@^��jp4ܳL�<HB��$�~d��� 6Fv0����_iB���W��F�S�M���T��A�I�?X�����>�P^��p���Zn�K�- �-�g��&�	�wg��3����A�7�m]���P<�����8T�F>T��\��t`�V�C��)ρ^�v][q��{�J�L�S�����HƖ�m1_�=��mbwa=v���_����ӈ&���v���*"a���A`!�r��ET?͞hI 3�܈_w�+�[7�����T�
?�NM(0(�a�i9w�l���b��)�������$2�I(9�VJ�Az2O
������or��m-&�+X��T�h0^���vo_J�'�s��G��9ұ��o��CkjyN����b�w��d4�u��)��$�>n�Z�S���j�q��ĺ]tڐ	�&�(�����*u�4 ��V������o�yE�pA���٧i�v�f�X�@��U9���P�CO�W�ˇ����a�� ��_��8NO3�����z��CV�yOjI}���G١�㨏���H>%��"l��aCA:��b�k�{B�}��;�m��<�A�t�*�k����Z���o@�q��U�'EZJ\�����|��Q���|?KG=܂Y+y���	}Gh�syL�7ʚh�'7����J֡J.��8���fX}H��;Qa(a'�_��5*�Y�+Ϝ}�uD�g����m��<�.���k�"`�|W���I���lTTky�s	��ڋi�}��"%0���)To��3g��@
v劀�Q���У��@q`0*^�mZہ����M4��&::�AiC�
#�Ƹќx5��J���&_��u)bε�YYf�O�>�!��C�S��M����� K����$IAW�]ɶ`av��<m�o�:4N��v
um��0��ߦ%�J������Kw
��H{�t����Aٟk�X�[%񬹖��W��P�,'A�v�])@Uj8�!$�KL�e+9�T�#I}^d��<�3؛�'gds���kD��y7fo='���璞�.�؛��g���)C������WS���$k���V�?$��:��
�H��Pu��X	?\�9�m�0D����}AA8���\=�׾D�J���>;�y��um�hqTS�?��X����kH<������Ȑ�\���짽�r�oZ��e�Y�0_�Ya�<-<���D<�BJRE�Y j}eۼ��t���dn?e��>�aN6�}��'*&�b��W^�@��ͭ+������&��]s_Q�J�V�Yl:�d�̏����z�a�Y�F�J��Jo�>�l!L�\M�W�+��ˬ.�v��Ԃ,-ψn6�T�я���!��4<��%vx�W�J���^G��J���4;^�T'1Iyh��N��.1c�����mDF�2��G�uYlHo��� 0rV���B�]��<�;�g��)`v��q��`B�K��_Oi4=Ħ&�A�`��i����i��M@gNY�O?�'�4-�ZWEa��`����IW9�g�M����n��������@��nI��4�N-�L�=Nȋn[E߳�v������P�B/��1��;\�ix�i���-:�(��\�s�qZ
�z�;,¿.<ZS8�)�~�u��B����۶�C-�y]ZE��'M!m;�%U[u���y��\�;��W��`C%�Pr��
4�6~F�$�����J�Xx�^e�`mB��,W��Q"�����տ��iRH�j�q%v�A �>ۃ�SU�<�rYVoŧ��N�n�*��y;�QJe�z�V� QC4�l�lS�e�x�=�jR3��V:��v�=�en��w��1�d�\m�ؘDk�X!;� ��[0����	�� #���$��z�DS��6C�ea��M�J���ણU--5��;��Z?~��n��VB�\��&r�cN U�oPS6H���H�������m�#�㯸|Y��r�*v���m���p�s��K�\��G���_����3i1W$�AEJ*��N�i����%1|�B��.N@(��

*��W�y����ZTSZh��g�H�#%��وlN�������j���&I�I҅�M�@�Lw�=��H%�θ1��e�S#B�/ģ,b#�挲2����N?����d)�ȕ� 曖�侂`վ��+R��48�ҭ���|>�g̺@��F�e��q��a�˛7��iG�x�܏w E����dEdT���1V���	�۸1j$
��U\�hg��tb�y��N���k	����8�����2QU�k�̬{Eb�r`�a$�8�����v8��j<8�6���˽�Q�G��rG�p;���1����hП4�����)����Yu1H��d��0��.�#:���/�v>l�?�=�͘�
��ȟ��tuC��&�<���A/��y�hz~����
��&$|��t��VFO�J����՘WP�ϻ�V�t��n#}t1/5eҪ��z����|Ǵ��yY0�e��t�^�+�f��]��ew;��;��bƔW^lWp0�D�����P�P�Tv�F]�k�p�g|�*r� ��!�k9q�F�3�\�T��T�=�iܛD{q��\�߄"
L��7χ%Y"3�IǒlNPd?=���흨��x�QE��Du7:ji��S�s����d�p��X6�d�������`����Ls]��绋�8�%&~-�Z@��P4����4�͙�� }�"�,�]���Usׅ9e"����f���հ�2X���d�ٲ�`��S�f��*�fцu�{ty9��o5��߈�y��U70��ے/H�eC�D�����!���W5y���f��a�Rd�X�3�����o{�U?CB�Ⴥ���������е�xRЃb��9(�T����>���]��#$��� �����bz�Q��*�^�6���lhPO�2�A����sQh�x4lw=y�">�"1�k�?)�P:��1�\�ު¿�x(�p�ig�e�B-�J�?�~��
����h�+�X�!�ݱ�����G5��P����"�|1E��JS WJ�;!�,y�7�|Sw,`w$wk�!{� �w,��è���N5|䕪�k1�G��A��Զ�J�&�����>7I�J� ~Wy���毙rn��ұ��d�_��NF������لv ���<�9):��	����m���|����L(�}�P��	6��b��:��ڨ<�� �;�kO��Z~Umss^��� ��2�a��vr��w.���یt�h}�/�$1v���⏙X�YƝ��ġV���T�M	��Υ&W���_�|��|$).�G�'q\P�9LIĬ�������zn��� d���3���y���lZ��ZpS�pؽ�$��m<��-V�$��=�[��Den1D*.�K�k�.	��_�},@���}(���u4�NX§�L6�d�[�'p���$�L���ъH+���#~�O�"�FD�/f�	y-��-߄H����i#���34����{�E�)�"��Z!�x�N��W�,�gX؉��<n��P�� ���$پ�Ƅ�D2�>����h9把͕����r�c��e`L��̰I�2�i��QÛ��}E,ٵ�IO�t�[�˩��4��r�����
��c�|T��HQl���h"�`:3i�6[0gk˱��w�d���޼��"�w�����)�a�=�t0J�eI��XC��C� �u������Ͻ.��R@��?��LЀ`�9�- K� �k�|s�cW�*�!T9}���c�����kˡ�k�O'%О��KI���pp�]b�D��hk�8��RZ�@�F��r�RY��X^��V��'Bj��v��Z8�f �9��kN�N�g�=
��*voC,����;�72�멫! �Up�\��<G&	�5��Rv�k�|�`_�����B����L�:
Af��{ H�C����+5�Ʒ��t��_,�g@�F7{o��+��f��Z��̈́!�+L�\g�~^���Pا@�b82��Y���)��t�"�ɋ�}>d�w��"��mߘ�0�0("/:�u���P�t�Σ�#1Tr.-������^*������fޱ"T󦝯���	�b�����.z���&�*Z�M��SkQk���v�K�w%�W���+�\3J�Ó8���l���P�xU5l���8W�0�����6�C�+/���a]g.�	Dө+@�G�yL���H��@G��Ǥ�R{康17�e3aV
�q���⻍b*"]�%�7Z�yn�X��dՙ��D����G;;�M)=;33&z�ɶ����R(ą ���~Z6� p����1���U8!	i�o��=v(1����,�����0�����3�oo���t�=�A��W�0-z����5
0��Ai'���*6�T-��#vmy�a��
�N���V.y��vX2�m��*$�[Q���+G7 ���=R�?�q��[�����:�:e���ӫk7l|� +�8��XA@჆F�Ш�U��h��)���G��p\��Ou���)�ε_3���,C��9��ͅ�z��#�w�D���HG�O��¹B1�>�Ҭ #�Ö��*�1��gA��U*��v�0����SF0wzIz�Ӌ��ݡ�DA�
�Y,�?��-O`�Ts]�X�w�� N�*G|�� K!y��>��͓#�Yߤ�3~�n��	���+�iZ��$�AL:��(�v���b[���}.;C�HC�[݀[�jK��S�O��|w���w��0��.O*�#��{i���d�D/���<,G8?A�!��"���hWQ<�G7��{�É[�ʊ#1��=��92E��,qvYް�iB$1�!PY���d��%���i�g��?�X�� 0����A�^�;w�\�	d�sM���%4d����
�Y$��� ܖ_:��L��?�~�0S�_��	=P�/���L��-�@�|�J��߰���A�K;ŷ`�'��1;�\��R�.�褗���>;�Ciq=����{�W���i�D?�eg%�ͪW�Ft�єj����~+79�t�'�ȹ��O��~�%u.�8W�b�7��������[ݘ~�t��r~��l�OH�R��'��?F��yeSшI��Cm� �Nh�"**�抪��L;�Y�ŬVg7������K�A"?�Fc�KrGV)t�~���8)H�9� ���H�Rw10�_l��n�L��F�BѦ������~yCëj��Z��!���R�)o�L [���˫)C/��2�A�LAh���XTX�����1:w��� �H�<&KZ�'���OvqP����
�:8���:�/�z�.��p�7�����u���k��k�A�O���9O�tpqK�D�#0�v�Ttl�H6�n�y�1��qڵp-o%n"�^*���uVJ�?�wO�yi>�����##�)�������"�R���/�˸�^�複G����X�)�uvMH�?��]q~9������Q���Ì�y��8�m�z��\�cb�M���)��F��~��t��ļ�[Iű�6H$a����c�-:h�Yj�^:������	�;óس��J�;�<	���s�l�'�m���w��ٵ�Яɍ{��ի���?J|)����5Ȃ���'�/<�2�������/����b�D��4.�*NkB{i��f�b|_m���b��Z�b������R�|�)�n9�[x�?�GAc�$�LB/�m���h�]
�����!,�%�[�AC��UA��H�%��4�DF�E���3;9��9�5+'}H�DZ���A;U�Gu�u>�(���^Tu�p���V%���4�
U����?u5[�5k������p��$�L�D�Ѵ�M������o�?�gpM�4���{7 �� eR7�5d�pǁ�)�+=���rc��g:+v�N�.D�[^>�6L��e��<�\V������YC��Ea�[߿(����f���g�k{-ksw��<oC��d����'d���A�@C'cO�
�� ����P�L�-��qn��
�8�a|��`�� 4��������5��p�z��a}+��
~ � �d�22���aÜzD��оB׶�$�F�0!��7������82�C�¬H��b��u8˲�ˁ>��{��m$R)�1����T��O��S�mU���{�Ŀ���@�qk
�;�~�+�ŝp�6�H���4�]���@�wp��}t������V�a��	�t������Uas���ω�[��V���dA���b�.��R��:~�J���f'�O������za�"��c�� r��0���>GMJ��A*�Oɷ�XX�Y��u����6�^���P[��؅�/|i:���m0�^�������_��9�2Ej���X�P��*Ӯ�1sj;yq�:�H"���S"�b��^�\r�c���)=%! �Xz,k�5Iף�P��!l�d��$S��o���&{�e��)3L�
9���l@Er1ɅAΥ�b�J� �j;cO���0��V�� �M{�<K�zh�g8���ԙ��)�Up�{E�s��W �(�E��.���p.����p_X�U���q:>��h��nhU�G��u�<P����J|(#;��ɓq�tЋF8�36�`���l�P:%�W�"�*h��,�c�a��|�6`gU�����8�{�C�kOG�o��B�������Rb�ZWDs70�^I�4�`yĂ5;Y�͞+ʧ�2���0~F��3���O����PئGc�+�Ѿ�v��cIY�;O�����O��� zt\�"��(�G�l���F�B=��M�������TNt�\m��׀�Mmc��'??!#~��sS9�዇  ߶Rf��D
��g��^L��q�=4��y��UH̊߻ԯC���en_OMs'Q�c#�㐛e�}�\4�ا۬g�u� {��Nf\uH�����m��`{xF�%|���X��eSq|��w��0�'!����7��0d%c2��]��ٕ��s�x��u��Tn$��@�Vc �!�{�˼�L	4��L����읎^]���bu���.S����g
��M��W����{�[-������*�нf�&�P�T����	���;��q��X��a�l��/��Rb6b��4�*[ ,V�Yc�k�ɢb�4�X�"�?Yh;�3ͽ�j�|!7k����W�WS%�D�k	��ovNB��t�m�=!���-�(xp��	M������y�r=[F�0�zZ�e'�E*uD9���T���D��]���|\&��ì�Y�$]yK �y�����M)_rd���t<�@!��(�0��W��7��ɡ�7����	�Ya�2�[S��  N�ֶ�i���E�"H��%�u�<�ٿfֳ�D����7EZӨfX9W.5�ӚO�f�!�5����Z�Q���I�*���ːf�{k��TpQ2�y��G�����w���G���Wo��Ї��q�&�d-�t�
�y?O���9��j��(ك�@�X�iԓ�?�Px�}d��"ߥ�Y=�����<[�����{���G��0�Zm���}�w�I�=,2'�r�҆lR~���a��џh
d��;|�"�!�jj�[��i-R�?�Shp|(��x��0�1C�w\�FV<9�3$26�<^ �d7�b�(�m�)�d/� �T
B����0��~�~ň4#�1�c��N���*U���
m�s������?�C�2g��͸��9D@�R��$�6�C���qƺ�i�ٺ��I4	�Rp��3�Уx��Ҫ��;�sw��^��`��	���H�Q/��uz'Td<��mt��KA*GL{0��)�� ��
5l�
�u��O�wN��)z����V���~cLg�Y]vGk�0��s�7���ո�W��%<�{���Cj��h��C5G�3Y{&P��[ݓ�[A�����Yz���H6�^���Vu
/���c��KRwH�x�3���g+z���K�l�(,zy@2S0j̦�	 �WV��إj(Nfr*w��5A���i�}-�fs�6�9�[oq����,2Hh�i��ʫ�J�xI����`ǣK�S�ޜM�W�w҇x� �7���o��J)R�&���ܫ��&��r�Bꀝ�!S��6���`2(�1�`:�Dc_�p0�0�������߳���������l���	�g�W s%b�������b?AYić��n/�^�Ō�U1z��.7��I��GY̊��d�����B����N�mv���o�=��0����cI�&۶�2v�Z
��v0)�%1,��}��^�!D��D��e�������E>|v��t(��8�w��1]�))巐���Z�~yo/m�^��*r ÜyK�7��i� ���E�3ڬ*�F��<.>�K8=c�h>����+���N`�l�M#F��I�i�����.3q�hka�q�l#[��>}���(?Jl��SY�&��Ω$o�K�P���Pg	��E��	���~�v��^S���k8��R0���q�-�5��=���XvX~5HW�B�uE�h;�I-k�.XܪOP���Z�ɷ�~�nߵqQ^Q�����ً�F_�Y�~H��i��B��XC}�;S�1O���˧F5 ʙs����6�\Q���Ǖ5`,�c���|�U8��@7��؂ ���/5ϸ��Cc���{Új*=q��e�ϔD[fؑӸG�B�U���m���\*-�}!Nㄮ�e'Z9ݸm��ԉ����}|�w'��D�*���V��s��e=����xL&�����v&�fJ��q����A/��1�����K��)�S���p��c([NM3� �K2~�WꯨIϺ�5l�-�~�����P�p�R�\;�#�I�.l=T�7���E��N���"�$9~�)�ލ��c�F�6[�Ϣ��ݮ:�I��d]���#Z���K)�]�WA����F�,x;�[�'��1��ɛԑ���<D;�u�a ����B�����r�nTw� ��p�$�+x��8!ո\�����mYJ�4>iX�&�5˼5���>�D�j���,��9#O��~��)����tJ�`v�6�Y��\0��|�������=Gߊ'��F�Y�A)��uL���S�^�/��ɖ���,zos1����7�f�bj[��J9!�:7sx ���4�#&�1��1��׷h�]��Y/�j�(�c�^1A��.P��F@1���W-;L���#�CR�VڟM��DB�_-��q'KP}Ra�yY��k�9��m2�#d�0)v�W�i�Z�r�H�Us,Ђ�xV,;L��{~�d�J�p��Ya�F.�n2&Z*pˋ���9pV���<���_��ƃc��5S�ho#�`��r��/�#�6���px���X����_3.�r��m��z5����͹���T1��� v�L`O;Z�.8��.�WyϒF��� d��ڴ~U���]TT���[���OҔ����g�R����%8&�rB���y&�k��Mj����(?Mu�h�I��"?m4	���f`�̓�M�r�Wt)3�:E��'� �3�D��B#Z�Zo$�Ȁ0�sa���l����^(�3U���O`^�� �o���$��`�q�A�}��B��H&PƓ1@���:t}�O������t~��� ��h'+9	3���vV��*���}̝@���P��#�i�hJL��e�������<���������X���ό!#4��#��I`JiPn���WQJtFǜ%,�4���;R��;�_���1�>;M���'��+Y����0ϛ�?�]i9��6G�z���N��m�mRШ��١� �ah�?��u��$��կ�� �����OzS��s�
\@31HrĠ4}���.�1P����˂���T~ƅ�n�),����j9��-5����ͅ� ~�s8ef$�m[�v�BX���#�� �F��'����sQm&����أI	m���Uְv��y�%����&�SOb�
;%
�f����́<�?�"P�%�	$�����N�p��&������,�l,=1p�Z�3�?��ȚR>�d�P�I�XB�Ev���$�D3�s�n�W��k�I��za�ɱQk8o��f��6f���T�륦q����;�i� �<���`�Ϸg_E��B�1LK`�+�f__���]��V�h~�h���u�m�K�����2�z��z��wcJ�����%q[@�x%�ʈe���h�rd�D��	����x~y��u�B�26]W�Ƭ��1 !�I�gai�k��eg#&�K�=Ԁ�)�f2�*Vp��&G�F�T�%�c!�#q�9UCZg�f5Hh��g���vB�(i�O�ۈ0s��e�2�]���نʲ������s�cO�eh�P3�>v~GV�	��22切�KE/���]vL��]�_��-��sf�'�Z~�Ƃt�V7����J ռD�VX�W���^������ÿֽx�V��	����U/^�.y��6b������u�ހ4[	i�C�D��r��r��K2!!���{���Q`���Aָ9Bm�C����zWa1=|o�
/)�O�8�9�v�K���c�D���!�,�zv�-��T`�|����Fg�x�|da�F~����*�N}IW�#`O�b�r4ň��c5�/	�&�!kE��%Z�����If��?��۱t�;�)���-�i��U��-0��{�EG��rԑ�I즆������o���j�T`�"GcP����^�n�J�{Dh&kD��P�#��	0�b'� L�y�j%lW��������+G�7��p��h1���f�[PE�"q��cv��.X�ƛ년��,����%O�l,N랻�@sWX��Ӫ�6,w�sЇ�}�y���3�~yl�fZ
��F�`F��;K߱��>�e�D�
�:���U@gwK��j��ѹ�d|�/�M�٬RL?yd������S �*u��=��-��w�W�4@
���΄e�m�V�ȽP]����8��A��I� �ȴx�ݙ����ऀѶ�p��ծ�=tK�O��;ڼ
�0{.��Z�~��f�8C�I���)��YF�a�
�cmp�¸O~2���ܳ��6����F��};�]Mf�`4�R�z���v9�O����OV�c&�2A:�0�������-�2�I;]'a~Ա�QvJz�w����N������j��y���R���h��>=Uj����J�c�:��u���ת�޴l��$�Jk�fA�|�vM�PϮX�����#h�AC���6ÿ�M.�.���Z��Cxzq<��kH����}�4�L�x�Ff%ҟ7��b�:��?�k-��px���M>�]Ϛ1���d<�
��0,���y[ 7,�x�*V�vl��I���}~x_U3i�[��Q.ӳ����M�xAp�xN�����ɉ��
Ov��P��"zí���h/b�AtM�v�Y�w�����j&� �tK���y��1~��\,�&���>��(z:�j
�~��F��WkdWtHS2�͸ѹ��|�}�%�<����+҈�F�X|cr=�JX�3	���%�5����������QY��.I$T�}��CE\����mA4�����B7z3�d����n�=^���F�}.����y��x�6"u��R┸8�y�Zޭ��	�$�Y�v	޻��&����P�[/s��2�&HE��,��>���LA8\�w+`�
2 ���}����e�H[u���jR�<,a)6I��6�"�&�.A�Y��\��.��>���`\[��k�{�y,���J��ـ�����ES_d<����w^m7�n� nj9��<���^
-ʥRl��A'����b�`���7"�(�4�5�����sDbL��>��͋���aW�
�-�sCE�r���X:\À���� w~���Oc^�N L���[�p�a���"���kզWbb,(yp_nT@��64ӆY����Y�,mz�kSβh���?�
?�b\(�ak�R5�#0o�՘6��|_O�k��W�G�-����������HH�*�/�ytD��>2��w����8F�hG�=�1b5�a��/�+3�c�'���~�~���ܧ����meh�5ߪ�Q-���5���a�d��!��W3�l��F�&���6��G�&G�B��ᳩC��g) ��[K`.aڙAlЕ���~	�*�a�+�:z�ё+�8W�����?�L�l�U��
��S�5ȍB���:I"���I�G��Dd��,�x4��f�z��R��9�
Ca���j"S";K>z����������t�>B����0)�/�n�O�4Y��~�3����`�����9��SR]H�c�)��35��B&���윉���vDB{�3�pXF���Xm)�M��K;dH��<Q+u�"g��y@eXg�Ĥ�#��j�x����wڌ*���k1�������DƛkĹ-:�Dk���䌟9$x<~=&���)�ͳ��I6��CT�Z��/�Z�87֬�6g�|��``6����`%���]�KU^���<:���/�3�{%W�j��4���pVw��Uނ3fj �/�l�fe��+�;Ύ����*@�2A�-�4ظ��B�a`0�8nܛ��s��?kY�E��kq�kd���F�3����z�	�;A?p� ����?�z�x�KKJd���JY%�SBÓ����	����C�>��t���sLo���Mf,�����i��[؁ɛ���B7������pp�����L�)���1�mAT���Q�6v�x�<	��=p��͢#�?�Mp�<W �Ӟ�WL��K�t5��J�:��'�Op��"���0��\P�i�ㄒ�ę:�l51�J��1�V	`��&������.˥M��I{ ��p��Qᘭ{�����:�s�c�&��Q`�"SX���j�T��\gI �B�a^��[�-���wB(�Dj���x�����oBY�'��y̘za���<���W4��n�ywD�il��C��ts,�r�ԙ�(PY|��>X�{e7��/�oX^�Gc�O_�x��>����S�5$JB=l�A��;,қ��
�4�R?UP�����ײ$����z	��9�*j�;�i��D��݂�W��<�0���4r;uYm@!d�ޝ�F�AvJM�ys*�d.i�t���#�@^uT`/8�K�d����s�Zk<�š�@�~\b͡\g+ld�s������a�n�x���_q �&�����Q��~�W��SMƮ�4	R`�wr��.L���W�$I�#	>�!K�M���`��o��_�,�p���˩���m�Ձ�2��Y�F�5|hɈ�$�8I@
�,��M���6RB�I�߿�Zb[x��V?2lBMw���>&�9�3E}[�&Ε<"��쨐_Fe��v?Z��:D,�طME�֯~N�J��iK<�xXz|`;>����@��r�F~U��.6u��(H��EU?�'�@!�+�.��P��O�dJL:����ijUm�0ԓiK�>�Ց�(�Q�mCq�C�����Z/׬��&�U�EF����2���Ŗ�Uн�/.�ҙ�F��:m�Mx�Y�f���<�n�����#�P��_a�ǚ�9���?�^gg��j�>���=��(�����Iw{b���(Y�`@ֳ^>P�|$�!x�;F-s騩�Y��iT�Sm[�3Hƒ�\sJ|��[�嘧�n��H8w��(b���M9��3V������-8�ʔ��(3<f�ID& 7~^X��i��`K�/��KqL��%E�{%���w3c�v�PsP����[����H}��},�k{��jmD8@�~�*���fd�7��q������{<�*��5��Z��}�4��7+l��-����;�����v1�KX7Q�N���q}I3`�f'"�{�r��>K?B��#a�g]�s]F.�*�-����샴������R6��Qֲ�s��_�(�*�n�Y���oM��J�pO,�������
�e�u�*�>�ؙ@T�;���m��P�v��כ�xߔQ�2�%��jĲ��aAVQUJ�V8��]�O�zG5�p��7��$]u|�(�Z~��%�7���^�����$dG�W]rm����W��]���G��#�D�x�#N��qd~i����[���d���6���3���-����,z��9�+��g�a�3a/�4xjlɓ��Ef��/�B�@�G�%!Ȍ/͸e�fí�8���#��֨��>�.�~�Lh����w#K�����h����vΏ߾!��q�\�i�*�WR"C�p��&F��c���^�<�1�#�M���0[녲��O_g������ �ȟ�<=tl�����ǹ,�݂i�)��Tm}�x�_�ҳ�+}�|^��*�3֪h�&��;��7����T��<+-���H!�=7�:������k𶧰�Y��ZH��X����U-ʭ��v������B�~1h�bP[�n�h���E<9���%�>w�J� ��3S	}�D�5G�������u�Ѫ����s�A|��F�8fh�`�1V�k�X�w��/��5�#�3�xu&���ۺ��u�Ԃu�F�7�a�T��?���?��)&�Q����𙫍�k"U�A�a��m��h���L��~r5�a|����B�8<�Vҙ�qi}��F|�����D:�SK��)2�� Gs�o#��m	 ��ѹ�lŤɯd���보O�R-��;FM5�\]v���l;��,���
�y��x���.��Ǟ.4�N��`&�5��Y&����m(4� �����Ҕj��\���Ki����ĭ��K@u��P��f�7� =� H���+�J��h��<_��f�[�Vf��=��Z��~�'9�u4��#�~���!�y����L���6��|���?S��4��	�˵�J���L�=9mNw����*$���N�C�ºtwߙ��C����ϔ��ϼ�8����^ԛꘁ�s��MJ� &25B��_��1��3T���[���ED�\
>��O�oK>���8�(�ԛ�4ٍO����/(h�	�X}��^�D����oP��h�>�%����)�#�;���I"���ﷳQ��!Bm��T�R�	�=����/����r����/�$]H%'���8.A;��U~����CȐ���8|i3A���x">#y{�٨��G���	_h��GJBȟV��t*��}W)��L�P%˘N���$fv@[-�LCΗO��zv�3�����ʉ�?Ϡ�A'�u���1x���v;n�y��X��TR3 ��LTh�!��&���p,!��쑓�i�*�ͼQ߾�C��3�X��+}w��8����0�0�ii^"����qK�aw���(y��$J�Ʃ	� ���.*�?��䀅��מh�k�����5�x�W��C��O\�!Q0�z�V����*=�]r�6W-L؞+o�o�.��xU3��[h��wIWS��o�W�)占�k?�0, �=a+6q5�ƹ��1	V���n}8� !S&� �!1;�Nhr_�ƥ�쬎N�bI�~�PX
7�=��h��+�uu�J���;�a�e���56�R�H�:S(�(���Z��)�?�Z�¿���a�k�E%l$�Q+�0�r�@�}f��}Y�o>�8�i����E��%�$G'1���d"C���Cm����`�
<���3a�ՑJ~CK1�c��g� �;F�(�uԒ)�9r��+�������J/��·(My�/T���Ȩ �u� �t_쯓��j���B\�e�,M���q�ⱁ��hk]~�ȦG����K?=V�f��"ϐ�W�5��<c�k�l#]�f��^<F8A�
�6�r�7\�
�3?,�; %�M�kŖ��Pڵ>����b�y�-�2tc��}���O�_���F���<
��Q݀e��7��ň讑� �;�c�t�x"��))����a��[2����t��lؒ+16�'�����F���9��f�MP���L�}_@�K��%/!�Rq.'ѧm~I��>I_s
��[�=��V� (�&5�Ye� ��m�5v�W,u��C`Ϫ(r}�}�Ƽ�cɻ���������i�[�j�Q�@��ET�����0��$�f�6����B�,����22�)?�"n;����@DC!Rd����h#�@+����f��GS���OGŝ���P&��};nx��b�:��A��o��5�9�tE�f2P'K�/i� ��9���a��g���q��TF"��Gq��%?�#E|.O������=˥���T���X!�&��B��"'9.� ����n*�O��qA�Y
��gg:kQ2����}*��Yh�2Kz���r�zM�^�wX�q�\M7x/?h�����_�&�nl�f?�ˉ�B�A�l%����"����y8��%��7j��@Wҙ��TX^<�ʢԛ�_���Ѳ̏�Ä�Nߖy40��V�t�Skd?wobj�I�S}�i���Kh���eH��0V����1pjp�� '��*�?�1��:�)3���!���y1�ϲ�	ll[JI-Ɩ)0%�z��
���i2ĭ$����ã ,�|��kD�W5�D�o! �ȞT2P�`׾8�øH�B��9)������>|EN����2~�G��T��̖��]_�}g\9�V�G����\���$3��$�_�Y
zL=.��h[S����w�&eJ���R�K��Ȥ��ӧ�||�yd��B;5��|�X�T;R���t�5� �?"������8�H��g1^�ї��{��s�_�2tl�rA�ݩ{2:��XZq�^ۨn�����/� 홿]�+�:���Z�M3�ק��^P$	�nz]?��{�^��=��7
�Y��|@焵hG���
�F>j�)��� \
�7%%�+p&daZ	�Wü9h�	��v�B�Qwԛ���y9��i|&{S��:F�C�E]�j�M���J�`{'�!&�3�6�Pjt&�x�hN�py<��v�4��=��d��Һz�~�jf$��
���D	���4�4����%��K�c�n��7ff��YP�_�����(�����>����h�l���7qp�|�־+ j��/	2����)a��%��t�!��<щ�9X�+�*s�#T!�k�Ny���,)7![���S�,^Wq��l�RrYqڟi�-��bJ+��9I�D7̕M�gl�%7����#o�/��P��<%sЙ����`�Q__��#���w����X�嘖$��c���<g�M�/��R*?�ݢtF=�g5�ߡ�n����A4c�VO�I�Gݴ�}j��w��-ܠ��S7�^Y�Ew#~I����%�Pn㼛YrQ�� =�����1���:�<��'s���'A����A�iH�JI��v7Q�SHW{��y���4��O�mc��Q�-�ǬhPv��Q�/+gµ�#�E����7B�jh�c�}�\\f�!��E$�Pj�|#j�ȯ�ݜ!Wen����~,�dҵ6޹�S_[��1�F#{�Pb)	�z}�����L/��t~̡��"��]���p���Ʒ�#U�g�OMy���)�py4�����0G�K����i
ఄWj�5,m{rzv�1T���YE���~��1;�,�֒i���jO����b��F��0�+7��qh,r�D����=��)�S�y�����1�.��Te�f�RO/jy�N]<&�29/C?f]ҳ�����"§$��%�٘��N��j0��Ȫ����!V=�-V�4�X�h�����w�!��N���ީ�����M���#tp��d������_�v�嗝��nI0���]�c4狙��0��L˙KBKq�A�e��f|E�\ꐢy~�a����x���+�2N�i��"%��B�W�����t��mY���S]+�nn��1䂷/Jǜ�`�����b�V��/�I4B9�bA�8@R��|��a8�a��'$�B�=�W9�s��>�a��V����T��D9x@�߻���Y�đ�K���-ur�������x8)	>�\M���B����fw��~(�\�8,���I��F�f��Z�.�s�k	�N�H���5���˪�CN8��5?6(�������I�t�'_tn�Dm�;�\b��f̅�8����Wp�U�X�W���&ײu�)��8����DM��<���t*�kv��QR�1�X�b�ݳ<ev��-����O'!�[�0���?�1O3�Y����UqZ1Njl�X �Ѿ�˹	:���ޤ3o�m�$�t�zn۝`�_��a�}Of�J_�4{�{A:o>�O�l�>E��l
���W4�D҈�����^�3_+}?ʝ&��񠒷�ő>�w��N�^�Q�)	���ƐB"h���w�>+"���`h,t:DZyJs��p�iE㜔�Wu��X)n�X�j8%�c�. �+RҴuL�b�>�J_�kHz-ZN1�f�A/Ι�OT��Ï����@����^F�S�o	�<s�~TGDe�6���/�63E�Eگ�C-��%zl (�1Wj��&
,�Oz��u���<��ގ�:��ѯ���
�;��,:-�՝�qS��g�b�/�ö[��X����w: _����B]62{���ر�`�\h��?�exI��g�$ �G]F��pⱭ��~�u�m��|��_�:���4G�'�H|����P,��G3
��9]����{� �XX?�\p0$J���n= Ԗ����@��u�A�b��&~y�=���$�4B�~a�|��PmA.��A䋯wһJ�޻��f`�t�q\&��L �����P��)�o]�Lڢǋ�w/�mΑ�c|�Sq1��v?a���"0��$���#��ʝ� ݎD-T��Ԑ�v�n=O�}��J������`+Y��K��� H�H:s�T��.9��.M'��9ZŬ
�4�:s!d�['��c]��Z~zi�e/e����͈�{�(�t=��_�l�	�k(�Ύ�kq���e��ݥ���fm��~�nz��<���Y��J��ؽ3�;���n���.
?��!\�,���)��a>�W�Z��s����q�n����N�zL�h� ��%�<f��l�
��t��fej�FE��:�Mt�H�����Ƕ��!���Pm\K���l�bQ�;Q�S��fE=F�_3�<ƌ�N��Z�ZI�9i�$�����{7�y�����W-�Y�ilBiD������p�?d}�����g�� ����J{y��m�&��]$��!T��ի�k;m�2V�|�ђ=�`FG��A��6> ٝ�u�����l���lƒ��? �,�e~��m�T:)p�Y�7n�z�oo�@?�*u֩�cң��2�h� `�j��Mk�3��I�K#�?KZ�{�ap�'�{���+�f3v��U��M����޷�,ܿ�v�Z�y� ��m��7��7���A��8���E�V!��eYx(}CŬ������{����^��E��J����-�z<0�����#��z�p9��_$�䞘M4���}��|�s��!Y�p�1�Aѧ����GN���eo� ��{�U���sm���?�s�wm>ʓ����p)z�e�l'J�*�O� �}u�Х��Q���{wq�T�1���ǧ���o�������1W.i��BIb�����X)W/tp�C��7�~u82�r��bJ��7��|^�s0�[ѓ��7a���n�])or�~��\�繆�˾X�x��ؚɏLM�ް��.Ó����=�n�'���OX��&�b�u������N7G��3z~c�P���N�#p�x�d=ݫr%<�X��=��ٔ^����}�z���d;eF���=�i{֬��;0������៎�!R"�P��R�e��6����<�,=#奱�Tl��iJur�e�μ[*�����'n���0{')t�/�Z ��"<��Db�E�����׉�����~�Ơ���
��UX���@3r�	���t�,R@�נ]?s̬ڋ�	y �R�zೂ׈�@���w�*��`3�'w���w
p�¯�}w�Q
j��=x���9�����f8�^�ȏ�:�,7BnU�-����/	���
�[����XL6����m�7��1|��l�XzrV?��]��&�������Jl�=K��;y"=\���bH�!�kJpP`���XJ�Es��Ef��I?���n�)$Ό#D�7�и��kq�� VQe�Xĭ��[ߦu�U��d\E��_ji;����jr�b~��B�B5�Mܙw��\�o�.���@��ئ�g���RyÒ�*f�Գ���T�i��!�3:�֚~�W߈#�b�'`��+�e�-�5�)�d�m,qg�g�>G��S��bT�6h,h�_���+���F����h��z���Ȟ�sV�A�ZZ��s��T�_��4��H�i���\��t��z�b0��o�'z?q��
�`�e�I�n��!lq9�8	`�B?���2J�0㪺G������М9�x��]��1�>&]B��Z%,�(pe��`��3��!��H��?�� ���o�Mt�lK��m�D$��?<�xPR����@Dl��g���Q�6-�;[%������7�5g6O{�"���	d��-8?��p=`����r85�,�s$s5��s��ճ� ��z���x�\ �M~ݰ�w{�����
0�������h��$�NW}N���#��u�&��|
ŮB ����B�щ���I�+i���Ɠ�x�f�m���HQ�b�m�-��w8Tzg��{��g�a��a�ƬV��&_��+A3�/�������ֲ��E��-"��@�:$�?�1bo^���!�C��;ofd�i��,B��Yt޴���\������Y�_AC�\�Z,�:������e�<V �L.��Y�tdF�TGL����e|:v˺�C!��Hg�J �~���S�Y'a	=�1��>T4'�WtP)+1`��������� @�yM\�q�
ƍ��3�ϾAH��������]��,ŨJe��W�ft�}�2+�W��ڹ���F(�G~��F��s<�_ns� h�굋G�ϻ�U;��	�����o9�̮���A*.L�?�=L�\K����폷ux���e���r=��ƞ���g���Yv��8�d|diiI��'Ī��9�q���
��.�<II~=�tf��5���(����
�Z/>"�r�X�$~c��i���r�tY�Ѯ4��"+�ւ��+�Uv�������n�X�9�����A5�ʬ ���Dg������)s��F���t.F���$1@�>�/hA�6�O�~P	�({�YZ8�(XAv����f�n���$0e�))�RQ��u��=]Ir�;����sJ1��g���-O��F��{Y��_~E�,+bt>������4��Yv�H�����M�ķN�r6R9?JqD�y�o���%���V�-�,|wt�q�E�p���c����lr�8E♵/~M !�1�M�^�ߠ��80�b	���{{ħ3���U%��)�w��uT
r#+^��_�'�Z$:��Ӯ_�X8�_��A->�H5��쎖	�&x�S�O��D�Z+5��؉Ʋ\����@X'��Ѭ]N=�pB���Rڠ���5�%��EE�J�����.K*�o�A@h�C� �X����	�V�`�&�*�ll�0����~�ғ0�2wA���ze�;�X%b[�5���/�\��GA���4�^�؂�x}��T����z6��x���*�e!�3m��eH����:Qig���;-m¤|�+��Q�Ųp>X6��ڠ�A<}7���a�5$�F��8Tr�;��P�E*s�e��|�Q`��N�Т��
�<����(�Utc(�չ��o���$@u������O�$��P��8������uQO�nX����p_�jt��g;m��{�������%��A�������J�wyڝ�~�j34ӣ��D��:p/��}觉��6�hw2� ��.����5tD��(r&I�\���ks�h2�\����̷D]^ �=*�8S�ݾ�����>n��7�'�H
:�/�)K/�(���_^��RP��S��v}�$Z;~H�U�B�+�i����uD�c@y��:: �����m�^�<�c��8�T4�s���ҵC�O�UP�N�>�k{x	��HtD�b�Y�޳�#�d���؄2�J%a(M4�Y�j����z��X��G��B�1:�|�C��z�X��6��""�{�-�!�D�`ٷ|�L�bwڮ.#��TA���e�0�H�O*�'<����퉾�U�c�O���+���U�ȸ��t���U}��.RX�B�Ź�DF���j<�sf���Ǻ	v�v"�1�-�l���.fcz|}�"�w���&�uic?FDs|ȳ�O�vV��8lh�gXJ�0BvÐπ�g}�$Ϲ���4�-&�0�;)�0��������P���ޘ�l��^
Y���μ��1^@��_'`}�Q��F`x;<v�D~�L���a��h�A����^�~�< ?G���D�;�.�sB�����&�՗�-�� ��I���M�۱�����K'��al� S+H��[���~��rsx����r7f�o����Q5� o��vm����*tI�E
���/�}Ώw���х,j]cX^U��4v{��jz=0v�l�òN���1Fib���+'Emކ�>Ā�@�h�����?����f^����Á��r��zW���
�)�uC�Ё�U��Ǟt�\�X5�=N<��L�b}
�0Fw�vJ	M�c�(K@t�Q�����8�o2�9���
ꣿKPiW�-W���2��a�ĭ���5�4�u�"G�d�g�)��nb�V]g���m�\eI�z!}J� Z�ӓ_�Y��昜	���P�;��I�F��8��I��׶mo.Gxk�V,im�`��Hؓ�T����"������']�s�?�nx��GB�^	�B	é��I�0HO&%=>�E��Y�����Y(Nb3��%�!����\0}�ݬ]�4����\��!��Q���O<+�h�Cˎ�4%��F5(y�2���9E�$E0��J�<�zuy��/Dgi�qr����̛�1Ɉ�/J]�UK�P@^1��MƂ@?���8J�b�hRr��m�� ��'��4��^K%z|׺�]!���X�:�N��+k����۝��t�'�'"J��9�\��u��w�4/wo�K��)�������yz|��y=&�nLV(9ȟi�_�.���]�"��Z�#g ����j��[j�K��F"St���Lo�ӯ�T�}�@�4�ԅ��<�̀�YLmV�ɚ�s�$�rd�`\!^��&��9��KW��ԟsӵӠ�l�	�ߌ�?�� ;�}�<^[^&��+Q��.��u��!&FH�L1@`0���.݅斐\�p�>��O���x�!-�=>�L�0��Z{�ij;Ih��!�I�;Q�hg_���O4#��L��Sp��@cJH�J���=�`�QUMʆ�U"��8�K��g��E���䳎Lb�ޡA�n�
ZF�������i��E1�j��QW#{-��h,j��Œͯ���Nu�Y>*ݯ����ǯ��A�&���#�1�\`����l��X��mc�pq����^�
���}g��&u�f����|b���iG�-/U�k��T�7�]}�-[�W��̬vx�-)v�p���2'1����4�� ���c�1�uz�px�=��pn�m�JK4�3����-<�1T���V��!�:�v	٥ki��2�i��$zr��q96�r���i;Cuf������,RPJ��a��Rn������� lP���R4�4UKsx��{�'�66:��,�|}opΨ;�`�6����]�07H��"���]�<��h�x����6PuM�u�1*�����N�ȇ�����V��v�l���f�֖f@D��C�~Ù@5~K&L�5xƢy}5�'h-�χ��\1rΒpO�RM���Y�mԷ� v��CXV���3JY�1����rכ���J2���-���c�r�#�A���L&Vr��Sj:aJ�3@ �2+�3��5��6�����sRϾF���M���ֻ
7o�(�`8?.���zzf��ԅFGÔtl�1���|o�4�e���_9n����gRŇʢ���p%���CQ��h�3��_��7gpȅ�@�����,(��K-+���a�]�:�D�QOr����1�8NoHY�a`W�.�,%��	��V9 ��|��NN{;/�7ei	nPQ&֗\��{��^�I�*�J����:�O�9��N�/�6�K
��i����ш)E�Ed/g>�pP�;��|qh����b{v ��e���`��wn�G�CO�ܭ�g�Q7}�R�螃���&Bpn�#���N)).NT���iì
&k�﬏E�e�R�Iu�-����s�#O��� ��FP�pO=]��'��]k/]쭕.�q��E����ZA:�S5�S{u��m#]$-݁7C�y�`�Ʀ�X���l����r:��9���[�d`j����6�%�P��S��_>�Cf�q���WTْ�	���C�ڵ�s�Av�"Pߺ�6޸l������������%��&�o�k������U�&~����s���ֳ<Y�qr�����dX_����D˅��[�K[�^hJ5�w<w�o4m�?KC�<�H�k܍x�P���{�'�s~B7�'|�����հֺ� \��E��a�!u�ߚB��w��۷[�v��6�m�Dgc�wHi(����&�I�\Q*�(~gq	k���{���8�]f��B}�-򦺃[���`�D��֖��l�qg�j[K���H�)Iݟw�U]�^<�M���"���$�I<$��doߋUkG*�	��c�w6�M��VL�y��\�^��%�Y�=�u�[�n�ti�j�ِ�rǌSf�*��&�"sѠ4ƿ�h�����^�2nih:+�][GX�<J�;���E�U6�;����;.��}}�������	�^0�"�@�/���p�x���{.�.RQ��G��p�KJ�b՞��
��k���CN�dZ
��mh��J$�^��I�-����Ւ��B�N7<Tq�F�$��oĜv�%G򗖯d�:PWz��!w4���!?󺓃�",��E7]J��`+t����O"�6b�"�~�ľY�ܽn�T|�r+�?�<�f�=xb���A m���m �������G$>���C_I����N}�������s$n�tֿ�&�7R�Y�J�*s(�Y�53kӖh�I��G��$o����8X��<(޿�z��ON�m//ŕ7\�M�+���^�KLݣ��px"	~nR�*]�p��Y��`·���]l}Z���!��T1��jϳ�[D��ӵtv�_�rS���0z耰��h�R��fi��t����N�6�M�|?�_��8�����l7=�N6m���-�d��h����-e���_U/іY��5/�fEr1�n��OW�U�9��,Lݫc�ǡ�q�\|�r�=���(Uf�P�� _|�FI?�!�v��1��2IwT�+��+�����̹D�ٷy; %3y�Ƙ�|�F�,�i��edO��"}��n+���ۑge��T���E
�����~����-����LNw�qϱu
fiW�.�"�e���'�Y^�l%�~�7�U���n·�k�����0�������B@3��V�8��������]�Q���-���5�BH�'���?�)�F�cm�؂��?�2����*�Zy�m�Nj��/0ZF_�^�ӱ5f�Mc���o�$��D
P��n�LA��F����y�N�|b���������M<㧀q������}?��#�J���=׵��#�����tQ���=!�J��e���S�����*.e��o��?N�Z�J�P� �Q½����֊���Q�˚�O���m	Xw6�\Rx��O.�\���,S�U�n#���;�_��k}(q:q�@�ۆG��.�C�Y�-�\	�ZOF��ż)�:0�ʭ�)�(�(�z��!yRf ��h��<������BZd��CPAc�H��Q���:'��0AZŭ��&W��K��\��
�v�Z�:h���	
������"?���
!���E�ܭ�I.<��#��Q�	�q����XdGĕ�`�	)��[�Z^�S��#A��4%'����7��O%�m=��D�o�v�K3��R(�H��g<w޽���"Z�v��U�*����Y�.f�Ŧ;䇑Z͋�W��\COֆb�j3�S]这��w6|�\�h�4:(q{nCv;.d�΢��&LHu�ʿ�,���r��.3=~�IOy�)}"(o������+Q	y��&�q*�`��b&�K�~"�J��Fs�u\*��=(�,:�i7�Љ��� �B��ȆS6q ����ָtX*�	������r@e4�m�l��ӱ�C��GW�"C�&��&,QW�^�;�\�����md	�����'�����텆�_X�%�Xp+n�I�'m}��nK���=�-���������P�L&���o�	&Q��qi3�d��G�܀�lYL���z%�`c$����S �QNx����!�_�_���טY��7-��d�dL�AZ{��WZ��.]�g8�T���Q���6��f�=�∓�^"b�4�ɾ�UUbX׺�O� $��8��>�S��s�{��y�����o�TS]A�g�Q��t�T5�~ ��rv�"5��+�(���[��N�[p_Ӆd
���D�$�[��8dT,���2��9��(�Mb��&r��7`��΂}��ە����}!{��B)��%�1O��Ru)�F���p����
�b��E���g�?� 0:.}���c�_���bZ�i�V�Or����_t�����
��S �SO�͂�������X�����ڞ�����+Wɧ����\��7�r.i��*�D�Tj�WNw��kIV͟E9c���0h�B��Gh�nxX��!�>&�%_���S�����i�� �T����$0^��2dH6�S�-m&�	I�0N �ˣ�|Aq�L���9���A�ț�xۼ��>W�1�	��})�d�<����Z@�MD��[MۏЛFϤ���2�[���ku�O+�8���dE}BM��~����g��� ��^t�	�f�6�����?������w�Zu~8��̋v��0�s�s�7�~��л���^�5�ٙ�Z����7���a}���GW�.߈�$�@m��+��k� Ь�&e�wNÈ!��k�'?¹&"�p�l�v���He��B�ѥ�/��V�a�;}�=bgY\+[k�Iv1A<�mF2}�3���_o����q�y�y�{�sƭ\��B̫�Mu�Z=
�v�i ��	ȘaC�YB x�ڏ�j���[K�K��qz�|�&cjexI�)}�i�M�b��R�cn���Cwt�X��Ӝy�Š���C�Zd�9c/���z	����(�,}q%����07�:�0�a�uq3f ����rd;���F����5�a��7����8��K�F)�N�3�����vq�a����u$ʴ*K��ȷ�Uk�ڬ~��5,��l{O���M����ٴb��wW��Њ�G+~`�<�`@��~�����Q��g����
\z腆�%���-�����@�c4k�0*���۷4%#�P������������D��T���&e�倜�x?�EU���3&o��7���7P�i��ˌ���r�P�@����D�(�v퐷����|W3(-�$�����d.Ƿ����NW-G�B�.;�"%X�e��9q����u=?�o(Ɵ/YG
/� *a7�9},��R�kD��e��h_��W�xILgmS#&F��V^n-�g���9u��k��Lot^�0���^�I`r38�6~*@���I��W�_�V�͒� �1g��B��_'n'�_��m!�����RMs�Xd��\WEQ( �������̡�[C/8�����J��v�^���4���\���=�w�n]u�R�w|Bb����"5�G�B�b2��e�ޭ�zI���X�Bf�Ur,bJ��]z�܈�֒�bZ����G���Ϫ�J$��)[f�XI?�U��*�/5?��YM�&���Kj`+ݘ�B~ �r� ��QFgǱc(~�۷�g]~�u�Y��9�Y��
B��7g�=�!?��Q6����:�GW��E�K!]uols{�v�X�B<��)t�r��1z��Vc��X�Ӷ�+������5zJ�[G|�&���ap� ey��������p�,"���Du�W�O/��1tS�&W��~�5 tZ���j U����]��̷��>�'�o�@� �jP�쒈9m�x4c6�Ұ��t��v6��6���<URQ�B����O����wnw���F`�4L�	��}?}�t��5.3n��&1���Q��]q7T�0tG}��VJS"��F2G(��w���J��rbW�	_w�e�7��uu�ݗ���<ɖ|AD�[u��}��9�+��a��+�ka]z�&3?��$B��ʰ��s��в2��Q�q�m�W	�[y�R��0�Z�r'` �\��pJ//�.ej�`K��z�h��ٺB�O��Ŷp�3�?h2a�_�K��z�L��;:�u��,�G�C����oٷ�+�����k驧�ո����T�Z�"nS�i�'��R���Z�NB����T�|s�)ƼY4�-�RE�%�㣔ć��^u1�o���d��r� �>��1?mt�j����I4��)׫t�X����"fv�^��VD�a��aεb��g�5�j5ٖ�K�Pk芿�N�*K��7]�]��o[ILY���K��1M�ْ7=qXe+4|�Ҝi?�̰
��lV��{?yp�.�^U�ڐ�j��N�č���D�}� ֕��� ���%�ݝ`Nu�6��#�]��"��kf��� l�����iI9Q ��Sb���ܲo9scns��-��K�ҫg�
6A�bkN�:\�M�5����Im������`�3}l4��H�&I�����}"�ti�8JI��J�?���U������*ٮnP1�uUP��"d��	��X5�iR�"C�D�����O5ݖ�>�M	�t�S4ԸB/�y[��B�R�~&c�ͭ�U�^�f:@ߌ��������o���I���8�����+�M�&Ãjy�]�i�̡�4���$�N
B�u&�����+�ﭟvi��9�t�u���6�1	Z��#Ä��b}�+j���C�h���AŇ�Qi���=���/��A�C�h�׉�x��vT!}}�-����۔q�;�Q��wnV޳J2�HLgd�pB
Ʈ^=0I�H�˜ԀR�5�� vh�+|���m�<��^a��?*�����v��֣��`4�i��+�Q)�����F�i'��h㺋�X�}͝�[�W �!��Ma�#Fy{���!�`9��1�Ő���U1U���OT�j���u�0"�5�dsϏB#DC�D]��l,W,��,YPd�:`����O�ߐ�4��[�V��H)�OцJƖ�l&:/���{�L 
����;�92P������%�N	a� F����M��� ̕r��:�n�g��G<͍4���}oy�Q�(՛ki6�v�����r!�';O
\�GFA��@�@v{/��6n�M���`��D�8?#_2��� �.��_�q����;��F[�q����'5֬͜�J��h*�y3�g"��	ڏ�=E0�v���*TE*�(�#m�����ԪD���cޚ��Ư��$��Ѿ�a_���2��3�5�H���J��!/�n��֐�׽/+�}�G�V�1$��V�8pv�K�fob�G2�\���A0hD�7;;n�4.+�r�q�Ln�p�6�����d(NT%��;��o���sz��+z%�<�ҴӹaQ9���ˢ�FK��0\�j�kïC�a2l(�nW����췬��$2�v+Mz����p���pLC����gf���kNK�}^���Z�	�ޣ���D��^�\R2�'��e�:r�����&��E�0���x�_�Ť,z0�Cɾש��Y���c*��G_��gA�Ys�F��4&�gC��<T��9��� we�G�c���|��r�f{��j�5jlí���"<���:~�-�'�˕�3b~�e���@��m��,��rt',��H{ �q�L�Yƿ��=2���&���Y�F~o�ɘJFڧ&���<���e'[fu�2���Op7d1�)��n'*�k����!�H&�.��D(��L��tn����p���x��pT5,͟�q�&Ϲ�����.nY�Y�K�i�<٢�9�3�/�>љ:{cL��5�P�*Saxl#�d�l���k��4{k d��� �9(,B�mN��k�u2��N� lY���:�Ԧl+������JM1.D��S&�+��7[-��̸�q��-p���AD"^^vQ,�>�xN����Ԝ�w%�MvλS���lX����C(�O�GJ��[��Ea�����إ#V ndΕryQ8-�/���L�����(��f�o�ƁS�үp&���;����9�!����G��Kd,`*}S�@?�\e�>�l=XJ��\��k��Zo��yws���ʹ�`w��I�q��:[Q�y�w��&G/ss��i�(.oj�!�\{�6�1B2^�'H=��n�:Am`�H䀅�!�2����
��l�o0<F3r<�!��q�V���r�o@��m�¹�X���+��-��dJ�^�TgSc 1NWZ��)>2ڒ��'3nD�Q^��L��`5-ʔ���/zFݶ�Ч����b�KUC��1ߊ�P����0B��#�!�`��"s��Iof�i~� �.��D���]m�Z>��<�;��^�����q��E�C�7���q���/�s�/
�	���߹B1�1���OCË��1��!��ʶ�1����l}����λ-�����({^AAL?�7g�"P#H�G�:����g�X}	#OP�!�fq�HD]��ǖ�S5>Q�a���T$�_`�V��sj y'���^H-�g~*�|�����N�h0|,'����gYݏ�7�&D�J���V=��&&����s74�; �`g8��56�kLPl�ե�6
𮩄7̟�e�ڸ͑�����V}9OC��k�~�Nh1��MHTP��ӮpE�,��,�y��ϥ�� �5#l�UӠ��O�������v�=F�D�Q\��(����Tnw���m��
�A�v�5�j�sRP�8K�? �\�b*�xY��#C �!����/��.ЕA}�
�x�/=���,�c��|ZX��ÜZ�Gp�u��޿.�������.Mf�9�D Q�)H�3ä�q)>�掠n~���_Շ�z�3WR=>�&4�JS�)��9�P������<��&��e�{7��?b$]̡�!������*��f��^�����E��fs	�+K/؋���q\$N�\U�+>{�,1`Gl-���b���rH����o(�P���a��㊛�ZX'[���PZ)Ou�Q@��
z�C�OP�ߴE�h�����R�M�"����q��j.P�?:�_�>qP��j-�-���J�Cy��*9>�N�{�����5���$�2c/K���iif9ޡ��)|��:��D8�Ǭ>��?��Y��ý�T3t�U�+L9�qQخkfI<m�c��"�#=A���j��cBf���ǽ����v�*E�Nܵ��"B��x�0We�
�����涖W���&p����%l�����]����N-��e�3�������&�
RA�%�fI����_���
�������i��bu��{*�0��@|��\v�n
ia��B��j�nI����v�f�@�]���P�z�
^�5֧�/���a�wp0�M�¦%���n��q���Nq�ps�����3�qI�3L�4.@{Ԥ�/9���QC�
B��N|2F�8���.A6�=k{I��9{�΢ X��c�v���d��1�oǋB-$�q,���a"ͳ��V`�
*��h՟\��$�Q��M��m��m:��`�Őt�K����R�@�8!�T��`|��vu��%�����b�gE�c4�b�)��nJ�1ì���I��]�_w�I�2�G0j��9�I٫�0�n�\�<��7������>./l�A�������I!X�O�P=�y��^��K�GU�IP>E����,����`�B@�(�Ĵ���f��x��Z�Ϗ����]�*]Ne� �e��Mb���h����`�D��$ 5�ǁ����tF[�j�e���>��0'P��ė`�zR̖:�������~xAFAJ\0 !=!���̶ջ�\�����fG�]���?���c?�8���:��/)��@8��b��=�V�l��:ʫF񨂼��G�Ѥ���چ�D"h���umT{t�K��g��h~l��b૘ب�|Ho�c��gA<�[�<��ދ٪�;��T�����vc1D�/^f�X��Q���qk�x,�"��sBl��������@��p�!&r+�d�S?u��P8����@�P�Wk]�1�)ؑ�Е��aA�cuq��m���v��6�&�X�B�|�]�zў�"�E�IZKk$ݠ�i�oκ�Y�v}�l�`�J�;ϝ�F��=�w5�孏���`Foݤ���L�o��X� Q����l��E�]��-�c���wr��Es�e?j؂ ���oz����a�I�<���.�wʩ��wKkޝ��oN�~V��E������p�5p��_h�I7sw;�ZU���yUR<���7�����m��bL>W�fW����_���{sD���4%�|��ɫK�s��YL��JBj����_Ms��[�1�\;�����O��D�n|NY��Nv�����h�|t��*ū`g0�Yi7���#;�W���z�8�L>e%$�{Q��@��B��Z��V,��kj�����+9�E!�R3�$-� R���ظ�y ��-�b�L�+B�!�WUZ ҧ^떌��x{r���Q�B������
6�	"�I�u_*�g/��j�-��n��~�)(����!��i�9)P$���<P�!ˑ]���qi�1&M�'���� 4���FVBja�"yC�P>��p�r��%��Y+�ӷ�������/�N��l����X�[�3��]�0Ҵ/��B>E ��DGz�^���t �r+� }�;�n*�r`��o+'��4�a�6���hx��{c��FҼ{��1,�at�=���jiWT+cZ����f$��z��0F�D]���%���"��J�L�`ٔAY���z����o{Ʈލ�u�|��F��(<���5�\[Jm���\��P
�SU�e�����[o���j��4�R�
T�ay������-���-�;W��:��X� ȁ����5��� �ij�㢳s�Jc0���!)���M��N��}њ��r"��?SY*�ܵ�S��%��Wh|a�g LC�r:�m�/�G%P�f*��D��c�R����@�`IO���5f�Y��.�_�z���#��� D��[����M�5"p�����ⷴ���1���OW�p�_��M��S�bBf�2�&7O&)ݣ�0�zCP��/˦ڤ�p��ìY�i��������oz�7C�v���Ikm�j�*���p��8�S�����J�(k0����ش�gdq�?܂�=���t�)�,�e�����p4)]�������� :z��]@��J�G$�:�.��/h1?�_Վ��s�����_�8��:�7x���k�r�o5��?�9:���fg��C�S $�c��- R�S7d�G/��x���Ă܌� ���;4�ɡ�"Y���v���\:52�֣L�>�	�mF���1/w�9��g;nh�6�6K=�E�2\���L;��~�?����
}AK�˽%K����E;A�^.�cɁg��`��Bz�a�h�¹�����bx	��ZW��ĭ)W��:-�I�����T�WRx�g�u�d��~��$P״�>Ί6�t�	�0.����_��M�,����a�STC6�Ƙ5ؖD�pcn 1��zg����-�SO���Q�~�$���j��n�m����1���W�\�.[���J�6�����Pi�!�����ٚ�UsY�9=����5���[��Ҳ����|&"��1�Aۯ�����W����M(�%rP�ӧj�cZ�qTD����WH��7�:�� ��h�������;ӿ�H1$1�a��4���o��g%Β#��P��1��ۤ��Sc�t���>'���a���Ͼ�Ò��iXyR-��t�9����9�uGo�)I�+�|��<���~��GV���|Q���v��f��Z	���]�m������*Ro�4�u=�H��4q� @#�B��ˡ�BҶF#������ܚ	���� pW:Q�����-f�bk�Q��) ~���5�L~<y)N>�l���"O_�e%�ŹM��d=��Ǩ�Gs�Y��(�t�%�;���JpQI-t�v��z���'�2TqR�gK�����@+*�!��z��g��\��IW7��h�����X��k����C�nё-x$��e�pIlGV�	�����6S5��,R3��W0u\�r��⡄���n�Ek�c([�SA6���J^o3B+�s�-�zP@Ct'�{�Fa���Q�XpM�3!�jP�����ʌ���0O�;w��p��R��I{�C_���{D/6}1f�(�N��-�����x͋�~�����Q��Y��W����_�$�\��7�H(�6y���ݓ#F>	Bpi,�ꔷ�m�=��;7n��מZ�|��ғ�5bґv�wH�V�75_��q�U�ˀ�DA�������������JAa\��>�qs��"�|J�sj_�X��zǜzg��Q��P�Que���9���!Î����[�_��8R���e���JEK?&n/�
�i6OH�4h�\r�֣+�H&��	�N�擠vi>-������+s\te��Hz?ƄQ��%�x�x.M���#:q�;Q�Swif��B�sIP��FF�"@�+͸�E��e�O�0��ڢ�s=m��b�F�l+B���.e������M�d�i���C��Ǵ�����{"���>���_2�.���9"��԰K���������x����VJ����&��[������G��L(��!br�#�L�6Ǆ��pq9~;Ѳ����C<  t�!�Ɂ!�����i)�+�2Zx�\��$ɟ���+�jA��^����OT4��"<��F�F�;沛��3:��/�����I��"6�L�gc��8��~�@��z�֖i-Xg5F�D��k�A)Һ��:l�q���}��(����m�\#}X���۫t�2���:#nqK��ŉ�A�P��A�7Hқ��"IgI��?�S��)��G
���8��s��WKZ�.�W���m4^�L��3h��]0�'/׀<�JC|�r�z\n��hrϤ��W!�1t:&�0p	;Xױ�:Vb}�B=�(�˖�������}U	3�F�xq=�Cԟ��)Jt>�<�ě:��M`2I���k��$b��qP�xsȌ����-�g�*|a�/N�12�)'Gҁ@�ϕ�~��h���0�T�Ƅ�kte�Q�h�T0@2�91�iU�hGx~�^	j�m�m؟��Bj����KM��;Ǘ�X�`��s�1e�uM ގ�eF�5�oof�z�[/Gζj
�n��~�jZ�-{e<s����z����l�4���"G�<�b���+<�b,^���Qj0f������C�^���Ԝ0��cu�B�O��Ԁs{d��/j��^#Ġ���z;��d�k#Ԉ�'5�^w>� ��Iw>�ei3�t��/�`CM3-�)[b;Nm�8��4s�Ǯ���o��Ət���cR�ݤ����r�#�ؤ��,����ȶu���%^_��4?Եv8�o�*�]��B��|^��C7���� ���[é�i�o��϶(��M������RP�{ܛU_�8�e�m�����z3?���N��ea�SJOep��������'�S�F�liO@sP�"܁\�osgP�j�R��e'ޡ�*d�t>Lǲ�]X��49u!|��p��u˽��̙�	(#-�8M����d����V�c��n���T5���_��~���9<DL�w���36X���q��wL��g��F�b6hg���S�(%8	вI�G�|��f맸gk݅"t �8B.P��R Wl�Imޠ�bq.�׉w�������I�NKY<3��7�`e�����զ_��4�4�JI���+ٶR�<�&�-9���!�T_z�6�q �F]��Tif��-�$j�56��8��R\Cu�Ә	،��H�»Ī|���LW>^́lɥ�pר�̃(��H�_4�"����?%BU��iaug�)/��	�xyD�f����:��}2�ȊPa��j�X;*� �A����iY��G�s`bQˊc-�m��*�|��c�[��.��a���Ø�y����*q�M\�[��ŧ4�XD��sQ�.���<N}���DbG7=�f7�GX����DӇ�����m��[��G��sr���W�����7��5ן�t�RUXxb�'�����YKN$]�I���n��wz��H�U�_��C!�<�#K�(���=-��ʜ�fys�K�Pv�w8��+���|����5��A�;,_g{�Pe����­	@ij���#�(-���X�Q�uU���C�[i�YH˳��73���ed��*�k���̪�����ٿ��0I��"�JGUi i�}�Wr\B0��逸�Ӽq��)�4�m��2�����L5:B��<˲ʾ��h���\�>�`b�da�	չ��w�9ӡCRzs�& !K5kª� ��%|_A('[Xu��C�:�r=�<#�{ؽ,ψ����Cɇ'�;WK%�P���Z���ٝ���=�*Bڪܖ��hH$��Z��DP�Km�u��4��F#�FӳK�r7��r6��|zY���@J�sl�������cw�ϟ���J�b
����DG��]�5s��PYL�2�����I��Su����<;���.�ePR�Б�����
"�A��xc�E��\,;�]��V���b��b�����AGul�y-C�O�B�"c��["k f�������i(�ݸ�8��4�+<��zl�D�+�YV�D5���+�n�]2�,���T���]i�ǃ��Z�t����q�����xl����b3��LDY�VJZ�F����Y{*�����|��)<����s�[s����s�9�G\�� L�N:�HV��^ƒ\�!��u-OTh���������nI*�,3�`�&�A���LN�N�=�ky�l� 5" h�,�]x�2.,���)���U�{�)�c�EϞ>�=�r����#[���( y� �va�A?�v[t!�B�|�����c�%Ѹ����O[��5P)��tM�[�91=�b[�����i��|���9\s�߷�?���F��ߔ�A��N��]�B�86���'S��V�UG��]$�+�!���F��Z%��E���5��b�~�C�%�)e�K�o��蹵�Q?8@�g��dٶ_~�H���Ȩ3��+��xR�Zn*<P}=@)�A��Y�;$!��W��`����[�r�鯖1����F �����k�"�m��$>�{�f�{>Wp�]���v2�����[�}q�B��y��y���px�4-90��SR.K\����2=ni���0�o����`���#�.{��8�/�r�W��<�*�{F�_Er	�G�If�z���Z��g�q,�`м�t�v�9ym!����bN%hc-��M0`j����k��,��s�W�V�օK�LH���%y)#�,�+Qϯ��\����8��;��m�<���ڹE��S���%�u�nS>q� &�JK�U�P��U�I�6Wn�ˎ� %17�/����Y��d9	��	��~��C�~��4.����m�����דd�������Z��O�D���ٹ$rM!滯A�\�y�Ʉ�M/�ח@r��!IF��v��.��RV�.��㠛���1���6�h��%��+	uwT%,�WQ#�l�-�e\#��82�H\>�(�;�`�w�Ʈ�:��h��J/�|��C�©������0���t$i1�g5���l7S�����Qj8g��)�ֺ��5��-��K7������9�������=}h�
������N �4�1˦������J)p�(=39}2}���S�T% �II���]+�����8�$�*Uj�j���W��0�f�df$�]�f��}_f]�gv��;�)��#�C���:���	g�,Z�&��sT��M6��Q�ly�H�ɟ���4mBm:�����sL|u�ZЇ{<�\%�"�9���M�(��b�RФ�/��Y� E����z��^m�Ǖ�L��^����	v;����w���5tC�ܱl�f�m���k :�VIrWh6���̻��H�k�W�8��ˀ�j�i�%����1��qy���*ˡ�inL����N��v�G4D9���������q��j�����������ХP@+B��W?q/Te�q ��;�$�s	2�$�@/¤�)q��S�_�9yS�� ���c�|'��e�pd�ڇ#g��2P�k��l-2%�V���I�C������j5�;T�eI�����"0 h�(H-X~��.� ��@ˊ\$��uP'`�����(�TD�Z-�gC�q(9�d�+�1u��A_�#Lym�2&��>b�$�󧞦�� ���{�<'/�g+���^�%�K�	�f�j����Vbw�:� �wإ�q�&�/�Ө�wV��[B�w躣u�����&��b@i��eN�Oɤ�zޝ���s ��R
��cc�-�nHO"(q��
xb��m�@DNO@,.�eMGA8AHYX�[�*�i5ws��L%=l�?��W�z:G�B-{�����?3'E�����0k����X��*���,䷪t)�%�́���՚gt	�.���)��T��=�T||���D��Nk�ů��rv`�����t���9��x���U�@�X(0K�3_�My���=��䛻��#_�~��#'���ƈ�:��C�F��d1dXO�P��ZvԲ�a�P���4t��Ő�����g��x��I��l1`�-R������N ^��V���j9�b�rv����h~�Kj�{��J&P'����\�D���
͊=(��F�"�R��������9���*�!�$gF�7u��fϺ$�2I��,�'��M!9��	�O�)�
��R]\��G.�)�.W�P}�
Bb*�5�z��B"�a�+_R�Ծ�x>ݒ�<��݌��n���Ҙ��k ܸ��9�7g�I��OrD�f3��V�������sa�Ǉ�O��1��3��� u!썮+'ͱ��ZR	�
2�Q�l(�پ��+J�)JT�*Ruj�r�o�I��Z��f�`G���,;s=���L��A_�im��70�$�mMN��~^rj�W�FY"m��
/�N�{����C��I��cH`�]ՉS�#�6�8��O@wRM��C~['~��m�������ͫ�Z���CM���I����X�W�(��P$S!֩SaJ7T�W4(Q.�R�s�Mpwz�y��qu�����;Kzrg-�+����p�\���8�F�t3�r]<��ҟ�����5� �	{R|�.l�����j{߈�*3� �(l�@��3��m�C>ռ-�@�[��Ű���㮷hc�FP�0倐N!� �Ԕ���~�&��
OJO� \G�U\.���1���ʖT���p�ܩ&��ĉ�e6ph(!���%˕�p�a��_�,8��_Uo��,�f�w���~��F[��#�K�(�s�O4Ύ�k�E��e;���H��1(�Z�0˝�b�����4"��	�Dmb2�U�M{� "{ �cp�%��'][��N�#L9�b�U���j��!��<�;+�5��lEk,�:h�B�pQ,5�&�'���ދ�,�"Å�J�kvM�h��m�']��L�(�5��S<`n��p/:AO��0��ߔ{�.�⡆mu��c�*����bE@Q��-��@;�|���$���2D��~�@r�V�]}//���d��@�M��dH�í�&D���1U��}�](�U2���ZEKu��L��A=m�;D]����j��ɭ� ���x��6�A����J�U��K q��Nr1���CS�6�%�x���yt��}�	C�_���Z�u�Z��&�Wo�0)�b�G=*��\�Uh�d2���f0�_���-�ąB�~(���u�g�,>q::��>�� ��^�X�\�&�M��Ns�H���$~��U��͓��D!�ۡ G���Nv4���d~]���.������"������U+g	5��넊>��)���y�&�A�V�T����S�]��[M������\�@Ԕ����gs��Miٜ݇�E4�
�&�Z�"7�/F�����o��8=��NWpA��
��hHF/���B_7���1WNp�S�o�i�r�e,��h��)�8�T�R�R����,��;�f t
q�g�_��Ƚ���Dv���=�^�J��65��
}�l���b)mS�(O����>�Ԏ��2 e;���i� �Y�������O���V(��_�է���.�����HHx��0��^������D��,�T$f���D��;��}ei&%lJ7&�<����:(\��B��G����-�iV#˵�����ڦ/��ǰ��f�y�����֮����2�c��:��^�b� �u����W�>rc��.Q�Ⱦ��)�\ʯ(	��j[��s�`�k�24�oVP��j(w��N�H��]�y,<+)N5%?W�����<g������4"�_g�L s�l��C�4
�^���������e����P�Y��5�p-琝+DRB��&�'%��+�١XMDZf�x<�� T�������bovry���K�e�O(g�@���p٥�S��-d*h�������Y�:�UI_�ٷcƷ���A絫��Ԏ[�J����6$�wgp�c�yq��`TYivX/�)�pr`�j�q�@��{$ )���qD凲&`uxg��bl�cm�Q���E���Sa�=K�ö0/��!l�^����E֥|�	��R�F����2�E{�߰��/�Ԙ�P���o�b�f��a�̇u#�$P��7��~�i�9
2�3�kD^mJ��+ s0:gB+����	c�$�`�+@<?��Ĺ�N��R�,�%��}N>���w�\�QEӕE g�/�ø!l*H��/�Z2��(U�k���d����	t*��V�mg�ЁB�_��*(�V��'��@Qe���03D��@W���^J�\]BdBZ���Rm:s�����9�jS�0���?��4-�_av1��?�ɐ��S��E3@V��W��Yo���{2�:�EGP&q͉��~^yٳK4�i�2��o^�Ee��i�9�@o�|g���һ%Hr^��c?'0G�D����y����]�x��#���5)0�.v�K��
+��X��	G�i#�'�A����w$0kf�p���4�������?һ ( V�:�g�i��g'���m)�~��cZ�Z0A/��O>ޱ�%t����R�Z͓*z�ʑ\&2�ɶ{)@�v�9$��?�ƹ�kε�'
�$���~�e|�A}r��}�������G*7��!�$�ń��!pP��(��q���w��8c���'�kSP�4ҵ=kFmç�P���A��f��@?�1 1w��\�y�̴֗���)��PPkw�9��Z�������?��*%�P��(�ya���'�t�!O�(�/xīG�ؼB��{g�T����H��m�h�ܱ���!�F�9��wN`�ږ�I���G=i�_��u�0*A|4�#�]����Wn ����إ~,���A��P��"	�b@kyYc�a�j aNR�	xy��5��S�F�"�<'];k��"���S%m�d�U?��X�A=%Tc0
ur� ��U�\���C�����A=�m�s�X�����# b�s��C ��������d�s�(����uI�k����~���Z������w(�^d�m�Npl�%"�y����oϠպU���8̞�#r,���vW��cSl���.#H.�؟{�;�]?j�~N�E�?�^���f�ޭgp��P�Ɩ��'��;_�d����$��b�l�"ɑy��R��vk8��*���?�y,;��?2��&t�Bă](�t��ge�#�Y����kU��a������4m�{q�h��W��YE�5�Hq��s� <@����,O�>��U�;��Y$�5�CT��i�n_�:=��&��GWA��:T���62f,Rәݨ�H�y�2r��0��:�㖜�!�JK#tp�a5�6�����XC���W���؉0��:]W�	�b����.�[�Yn��]t쟑	�0]o����V&4����/�GKa��rY��Z����>V�t��{��#S�6yC��1�o�Qd9��C�rU�?��8&=r�B��- �K������ڲ	qpu(�.�閄�p���:����H�:��yH�3%ߨ�{D��Ww���f8"���OM��_/Wv��x\�և�՟�] [��}!�1g��Y�3(�޿��C���� �q�>2}`�W���"��yOoι�S.NxΆE�/b�[O����c�*3��GT�;� '0���?(��B�s���VT���>:(P�9��]��W�*��YS���� /������8���~�P���䤰s��|�R1�BbeI�i�IMk_f�܃�>/�e��Q�|�B�Q)�m%�-!}� Sl��5h�2s/"Ҽ���~�v��� ���H�dX"�H"��,�A��3]�L�����ڂ&�v�i�Ξ<2��^��T�=1@�߀-l��,��5�~w�lc����G`��&���� �&���s�x�{A;��`��n�Q��g��M(�#�l�0|�\o�p!�3���g-饾���`��v"��ե�^������IdC��������@9��t�t���-������4c����&�*�̈j�Hk(��75�d�H�����Afx�T��fM�upC�8&ŋk����~F�,]�PL�MI5��=|A��3�t��+�2#Z��w�X��A&�Z�\{7��E�ƼBָ��ZB������������V�z�r�6�W�b�+G�.��Y�,�����Uԛ�GT�ɹB8�wn@9���\���d�P�d�	�/�?� 3UG�6ߗ��oC��Tv�nW�i�����80/�QKi
k}̭�����^��t���d����zd�� ��ٶ�'�?3��k��]�qxt�=Gh�h���gH���EPX|!��.�H;{���1/�/��U��-�I�K�̢��u2�k�����e�1el�xJ��<��Z�U����U�m����-,b� ��(��V�az)�?Z��CBP�Y^/���2�6��&խk�i"�����u�R�Kzm���2�qk�BW���Dy�-�1� ^�����������1��"�NWs�>��g��%L�,�}��#f� �ӂ��sw�R���P�q�r��6N��ܽ��D�-1Em4a�3U�����W~�f/�U�&�ۂ��D0߮�Jq`_��|��z��9gf�C�l.b�΀�-�+�6SS��*S�U�����t˚�=�=+��f��b��a�Lck�s�{��́��p�u�\mA�2��ق�Q�Zyv����E.X!��������e�=�o�pb�������5p��Õ���yn{eg��L���dj�=��I�k�8
SԠO����H�,��SM\U9\�fC������Us�2�'.�_�&$x�y�׭.��I��p�'�׀s��P�A���,����x��?����ܰ%��^A��V#��}粮��9��R��`���*
!�x���>��3�"~�o�|�4V�r�d�)�aW7o�4��ЎX5r���t���m��y���f]�1reYN�2V�2x��x�Ge�/�O�#pN\mF1�֎�'�ص�)��nw�9ѹw��3.)�\���9ז�B�!S�O X����o�MJ�"�w��ACj�M.�f�i��؃tB��]���<|.��:���n�B�ej�6��r� �4���G}�h�-D$���Q��QȚ��S譽\���C��lZ���` {[�W��7��D���� ͇��'�����j�?o�
�k��ɺ��@�[�7A��șA{�o�cv���뵐�$[{~!a^�:�����4��kl�A,E�����:[/����c����.��z�Ԛ0|]��D�|E6]�F��D���.�$L�f,��	��ؕ���{+'��ΰ�j���r����Mkw�aGƨ���<�(e������,�3���{�]�{�5��`�Y���G#��
��1lW)��Y��Lt��{��I$񇘾n4yp��p%x��$6i��Rc5��eP�¹!�f��:"3���|�L�ng-R% 
�
�;���i����,��pƷ�'���)��%pEW�&�V�ǼQ�L�L�R����M.xԲ��i�An�qt������?M6�B8t�CԈ��O��5{�e�}G��P}��J�V��X�QH�ZL��U�y�j�&��t9���K1��0�F�M�	N�zK��E�GjtQ�m�U~Ο���r�����6q�b3k�I����b��N؂���LD��>��.;�s%�3|���1Z��:��F3��}���ߑX��$��)W@>4|�~A6�]-LԶ�
#�,�E�{�F��^��J8COv�R ̅nE��V�D�	��?e��D�b����s��)Z<��,9��`��$.Jf���h��aG���M\.n�c;U&W>�,��0���,r�y�~�ϖ�b���E�;Sҁ��ޫ"���u�y�H��Ͼ9�Zs�m���jЩ.X쓃��L�]�H]j�_��N�
����
L�����إZk�|�`��Ur_ߣ�)E?������$�!)�@��/��d���5R��ْ��C�2�� �w��pI���~)��UP؎�?��O�L��\&vw��,S�bvz,���S,6f_��L]��]8a �����0D��:冨c��~Z�I�L6%z1B֠Jeq�Y�y�{�OP�o�n��[�7�W�~lb*��@�r7��V�(�Ii.�v�	h�N)��P�����!Z��lڰ�-�o���L�B�O,���Y�9MY8���~'�o�l{�li\�.����)�[�WG��9���gV~&pK�^�3�`k	'M�;��+����$���!�$�|�������D�T�7 ��1e%U�l�o�)y���+�]��ru�ertԆ�%|I����*�p`Y��ژ�Ɔf��L;(� �H�䰒���_� \�-�=�EpԱV-"D�K[l1�r�0�����X>����Ȑ|�q���9��G�^ �H3�_�2�&��0� x�,A������D�����筷����pLh��X-��8$��M��wJ�y��c�ah�"t���@��Ua5P^u{�]��(���=Y�MXk�g~��,�W��3����ki����P5�v���́;���%�%�uL���~���^�}���@^48�Pr�*=q7v�4��^@�B^TG#�qn�/�Ǻ�%���U,~��dc��)�fJ~{U������`7I8[�������2�F�"��J� j�3�Wi�u�Y��t\�Ze�볞���w�#Rs͋�>�%6��ȭ��]�4"v��� P��!>���/�{5�7R�3�A�<���$����(B.nLk�6��e���: �*]�hH�ucн���I��Z@d�x}��C���.U �J3��R��kD�6�����;��9ci����p=��Wa#(��f�!R"�����H��m?��}ɢS�^��?�}��KjO��x.������v�Ȍ�H_��,b�2>e�TU1V�ᐮbח�䒾���1dQ,PF�1پ���˻l�r8��0Ɉ&� g��Nl�؈vcڙ�X���ׁ%���ɚu��g���n�v~�)y�p������"H�gZ�WN�������{..[n�DC�UG�p���;�>���}�j�TE��SOx6�!$��e�3E�?���oMOg���<5�(,�	����\|�[|��N��P���������_�%�����uF�rH�^��~�X+E��jk�gӪH�V���Z��'G��0խ5�1��<d����h��!?��x�H<2�*6�nb�ph�^�����_��^n�&)�1^1�����n��tCճW�
4��EQ �`�_L+w�䝴��a�&׊��-��\5~@��\�g�|������lf�9��Eܐ����|�T2Z/��x��B+B)�h�̫����^���sr�.��U������t���C&��/����6JJ��.���)�2���<ŞB�;\=�k��>��ӿ� ��y��hd�d
��3�ݺo��\���ut�U��b�����C(��ge��n�!������@�&��O�imq��
�$;��&�h�]�{)Jx�q��/oAj=����A^I�oG�ٛ����t�KI�!p�p@D�o�F�1w,�PoMR:bG6y&q����� 9�kf�f[d�|gW�B��է-.Y�t�����]H���x��"@�(�#�����}���H~��++fxB�k���~�-y�ϋ�w��5c&��vs��`���7��v�A}*4$gʹpΞ:\��&vC�aGM@���Z�]ǽ�չ��[�t����������q��-�<���s���)m�ʫ�]|�k=i�1k��*&M�ž��'+�c������-g�PD �
zU����h3��.�T����z�5�uL��r�'����O�����:��U$9��L�f%�G�йb]t�u�	��i�GELx�i�, �%x�/Zp���o=K��w�+y���K�8�����V�vN?45i�^�dY�l������3p�*��x0\u�F�#0� ��*w>HcjS���l�&��#򺝕�6�Z��h�˵��%VGL��
�=�r���q��;Xy�v��g��[A2��\:k��)�)sC�R���9By�"VvY�;7`��K�=�ع�o":&�B%խ� %�sV�=粣�16y_)]�+T���1��AFx�?�Q֙���ߴتi�h�T���;p0����>��������zgPgFTԝ��{Z�&?F�U�2�������h�U7cxjǩ
��K�2�+�٪�J��@��[ؔ.?lZ�R�� ��@cF�S~�L.����Z�)0f�+���ov�:���SwFh\cE�(R�a��yhg��3��1��/����5�IOC�,cD�o�ւά ����4���F^��[m�@�]䓦t�p�ZOedv�U���>�O�At�4d�qiR�<�V��˱ox��T�Q�G^���t�#M�1��R�![��>�)�~�h� MU�f�d�oو]��a����]� ����A9�?�OO��̡ù���Q�B�B��}`�_�ۮ�)��Z��n�������a;U�v�Ѯ-��e� R_i�v5���u���x�u��|L�(�ōu�Fa|�.�C�/ﰤHuKfi�T����@ͿZE�����
=������8kM�[w�;#+�Ү�k��!�%���c�B�����㹭r�S ��O��?��p���9���י�(�s�vx�R��E�B�p�?E�*�灾.�x�{�� P=Bl��r��������*r�[2�
�=�QD���mdO�IN��D.�܍b�T��Sٿ�E��8����J����:�Xݓ�{��t�A�#�ASٜ���������U,3������^z=ԩ��5�i��>lL�2c�� �� ���ąg�)�34$�I^S�+ښ-�O��UBi����ƾ�3m���9��)>�Tӳ��Ğ�{%�
���y���tYĄ
��ߋBE$8��=G�?9_/�nw��Ա�˻#�;��G��Nc-�wx��0��Zj�x]7���g��t��x8�8������y�����0��fw��淂�2	�����9"���϶.R�k�3<1^�����f���.:-G�����C��.�����E�ըx��P;���6n��\�ER�aOt�n|�0��%D��L���2�i�^��T��jry#�!���<�x�� @�u����c#J�"�<Z[���x5�B���2b�,E�H�P�U�f�M��5�ګ$�5���Lp%�n�S[���]��s��؃�����Vp�`Z]�\��DLz}������q��>4���/�*�^r�l]z�����ŅQɍ�Mw�r6�䔪��#��xB�'�R�:�#U���V���Ú��בM��F��caӵ���YX����q�i�|���"_����x������U~��f+饝"~�ɦ�c-����=K����cF_beo��Y�{���^oD=�!
����]�j1(�V�����-�� �g�3���W}u�&1���t��������(��0x��չ�O`���6��3������ȧ�b߱a�B�o2��DP��2�̇�+��Q�� g�*.%34W/��*`;#xҳ1�Æm�|�{�� .�����(�'[���)	�*�/	J���`Iͅ�@��4�=)L;j� �H��@��}O�L�-��ttX��Þ�+@µ�������R� ��]pcO�V�Ƀ��{��޹ng�	�;�A�H�<�6�k�5��!	�ds{U��Ѕ�W%�(�agкh�Hqƛ8��sb5h&���Ȩ��e��z�D9�?Fe�"�����Qi��s�+-f>Pohڵ�������qY�Q����nը���4QW���3�A䣄#fzg�	��g�uw��5��2DB�.
v`r ��*�V��rX���M�~��&u���;-�G"�t��|\������� x�'`mY�E��Yn�4£
��8{K���\Bb1!~x~�#膺��]߀�y�t����߶p�����i�4���9��_���V q@87�����v��a����eI��fb
�;х�½H�9����!�E�������P~v3�w��)T��]Cc1$���ͳ�ӽ���Mg��':O�����瓐���f�����*�a��>M
�3���<ы�z�F�"~Z��t7S&AG�e�Rэ��uZ��.K+��]���z�o@�R�VGtg% �I��3]|�Ćɸ�3����R�J�lCc]���D��@�èsg=��q�n��pN!�F	�+cEg��x1�ۑ�$�CY5��'��}�|s�c��k]���ٿ�r2y�S�և̴�]�MT���{(�X���8L�����Z��*�$�X8N��gu:H�N9p�^�iX��]=|�Y��{#��v���@E����Ez{j��M��q��0]Nl�xV�B+�a�����M�'H4t��!� [��[I�à�Ș�f-#]u�� �Hl���z~���	���c�8�����#�<���X��Vs�Z�r��a6B[y �*���`ٹ��N�q�e[��ڽ�]����!�o��Њ���F8�˜���g�%��4�.n!���sW���}`'�+;V-��5���^5��bx;��\����G�DA$k��L�Sl�uрS����p�
K��0�	0y"x����ld��t�ŜL���:S���)pe;|�����葡���h=R1����:���2ed�8��p�U^9���֘Y"<���
�e 5�K�?W���5C�Pn>�X#����Ո���Ks
j`5MCL�_Am��Ȧ�晠��W�L���!��~�BhEs����+f���+
�KO�C�#�[��;1�d�)U���-L�&��{PD���l�_M�66�\B����n��/��Q�=L��]I,g��ߕA�yێ�ϴ�>X�����dĎ���bJeKv0�2�5���U0xv��h���"���ʛ~`��'����e�,.VA�+p������O�1P�#�^�䓇��"SS������1��d�5��P��(
�_5a�X+`K�����A6�m�0���'Y'����g���텃�]���a�0�S\R�0>o�����
=�-��*?y���MM��V�v/m2��x=�'o)oJ��6�ؼbn:�0��f��MR�7��S{IT �JFbwW������θXQT�q����I��:���-5�󛳑��@��%e"D�
^�fq��S����q�]d�lD�]�n	BB?��Ֆ�-�Q�g�#b��B�H�.��>�����U��l<��{rϮ&��{<�v�ab@#L��@s�, ��^�R�A�WUŠ���4n�~\mV���c0록���u��x�Q�BNq�o�����evMH��������}d~��L�%��sK�YcH���y妇�k�.&���k��N��;J%�5Mml�0��ʕj��s@��R�Y���q��~���Wy2m�B�?����;�贺;�QCwV�̕7�o��9�d�Th��gr�F|�h��k�>��L�/0N�e��2 _ϵ�ЅOK�͘��t��c߀���"L.$����&4!����G#�:Z�v�T�+� �"t���⥦�He����X+��ٔK�l���EТWf� D����ϱ�o�y_���ml�2�_����r����&�����M�����g��A"~`��ZUh�]�2�:�#��Ct(t��٩��E���{�4�M�ⲻɹbKK�$�1�b_b
:O����8�qW{N!S
d�tP&)+���$���C_D���J�/�v��sU�cٲ�AO��'�P")�:l�oe�|V��t�9��uhl{E�a�֦��g<[_���Z殖ۿ~q;( �e��uz�[
z�7zO���N"�MT��!�ɳ��1%Ԭ$G��c|(q'jQ%�x���x���ހ��[k>tμ��T
%Sm�t��+�Tխ����͹i����U�H�K�b�i��>q�	y�b��|9�Z�����(�5Ҩ��z'f2������1�C/�����W�P����{t\����SsA�m�i���8���ȼZo�ϧ�	LuB�er�I���
��F�meFk��	���}<5��j��Ú:K��GY�jFQ�~�_1�Ϳ�!�b?��p��}�2�$�[ө6���B�����*Y܂X��OcG_�<�>�x�VM�h�䶘.!����t�"�H�A��+�H٥�;ڃ�\��L��8��Ţ��{�.}�IΊ�>Pk�0E���H���͎>����F�)��`l���UM$-:�9�Ip�r��;�k�+�w�g�z����!�8����� ���g�/ff�q��SE�2c�ПZ�\H��
b"�K1f�2�I��B��b`Ѫ6�R؜j��=GE�.����j�Z&�+ƟUub�3���yh�|<xΰ������ lB���P��!�LfS��m8D��	��A%�u�]�#ڏ��t�r�J�b�1�b�}��-�u7nA�a
���7�/���s�[����vY�Ez����n��x��;c�d�kC-	�w�(�6+�کQ��\1ӫʮX�tF�@�,BH����V�wSX,�ȝ[F^��T(��� ���j;B!�(��d9^'sLl{r�=�=���q�5S^.�L�n�bF��+� H���V�_;3��燻#$���HAr��<��Fөk�H�[g�Z��Q���Ņ�~D��-���&R�Q_b�?�Y�6��HHH�e�(wl��ީwu���>�&R!+�+P�x�L��]������,ם@�H�g�Т����goA3ff/�F��@ˀL姹�u�Z��\,�D�_x��v`G%��6n!���<NI?��x���"��}�kNW\�!�9�?���N�a�/���B}?�o9"b!m�И��I=w u�C�h�_�I�T%4F��K�(%�RJ0�Zp5�4f�~�� �t4	X,�z�2[ ����+���^�	Tq
�>=[nJ:�g%TL0��/�Z?�_ޮ��DGu�썍%=��Y'pD�ɺe�5嬗U��jZ��� �d/���캬�*d�L}�$"uY�ř��U��s��K2�w�*�HMy�1Ą����#�n���Ѻ��#&�U-��/0�O�����`���b8l�N	G�;�p�fI3�ĥ2��H�6e2Gl�F�T�✆�;�D�w�Z�Dtxv������:��ճ%Bu��~w�T�@!�iF9��(��l�-8����� D���Gm|�2E��$��7�oa��Q6�&u\�L
�	��I@)\B��E�pa�,\p3M�I
*��+=bz遤�9���yC�,T�bc�!	�2��pYl�  F�ũ.�
�VV� �OhD�.���vKo���2MY�+�T$#Ϫ��1q��W"<�����#��s�rqt����o��U0���X��ǹ��K��zr[:�����0�K��_4�w"0�'������!g{�� @l���g�z�,
8�Np����#�Z�Μ M`�m�GP��w_vq�)tv@����5�&�Oθ��[{��$�V<��RG�!�'��wn����BvK}ȸ�C�s�3���˴���AӾ�Ǟ���0N�TnS�<��Z�s��L�r�{�j[j5ȵ�<��"ז��������:&�Q��Bg^i�9i�8m�Q�
3Q�ks�E��Z�-�љМ��QU��H��k퐜�Y��:`\������)5�=z��±��ik�H�Z�E����[��V�:�R�h�<&�Y�z�Y�MK��I����k�^9��_݅��Y�wj������6m���]�<��*��K��!�ڜgR��`!f��L��i���#gk�>�s���$���{��JMb� �3�^���0�]�:딦!R�颧ɨE&��'�
���1pM/�m�i�E�+]=�����!�a�K����i�XnSy��=����פ��ӫ�m�%�c�� =*[#�k�'����p����<�;��i�/��`��k6W)��m�U{ �`!�i�h���B(Xoxx�>�WQ��A'P5�ғ,N`�\@��sI �qoan�� �Jc[�a��B��w�@�aԞj�ݧ]�hzx��1���8ngUs��wJ"Y�/�xN�K�ڇXC�du��aeA�JJ������!�n�G�ʤ8HȮ���\��z��-���o�ܐ���J�1�����	j�����5]��jQD�X8�lc�k�˖� �����MH"L��p��"LoF�ȃ����2�����	���G�6o=�I�ҾԶX����������7.�g��^XsEڷ��q�8�*���˅�S*�v�/r`�_.)�,{������S��I΍(FK\mu��z��S�<u�$I��w�S�)'_!|��$0�`I��̈́��yY���ؙ��Ɇvx7x���v�p�m���ү���M:)��eћYc��+XE-�̟B���7���u'�E����V�(/˳�`hP�g��Wy�XMTH�7�iN�O���z��b"b���Ve폜KB��]���`N�T����R�v��ji��#�,3��:����g�t���	�8�~6x���}@E����|X2G� ڍ�G|�p����w}Z�'nsH�\��qTQjN�U$_��B9Ea9��-�/)��D����n{O����7�$R�=z�Nޭm��!/�w�'B�{��V����6�˯���;���(C%�]�DU!~���c��|���a|�������Q���ڜ{�t>{�D�F���,���QM���/��FM�&
��,��E��;�8���Ic}����{���5}�"h�D���N�1��A�Z�����'ī���<~�m�����%U��l;��Dz�m+�Gw\\с%y����/Ӹ��ُ48��a�|
l�P���I��G�?�7\��$$�%��Fs=�z��R�+S,���T��:���h?�i}W�1Ȏ��fŅ����J&�^
�+��U�'�����]�����iq���r�-�+�p���7�F�`�
.@�#���`�q�����n��u��b|�#�����cR�.X0�ӉK��W��	���dfΨW�S����I��*y������@���� h�Hd�1r�fJ��[�9�m��^�����L�Ü�r`�:#<#[�1m�k��LjKyُ�LEDLo�;��7. ��Âon&�< `�тñ�;o�m�h�Kq�ɮ�]��7(���9}ǔCn��&�N���}����ېV; ���k�!P���Fه'��R3�Hx1E��D�#�])�����RC�p\~T{*0��Ƃ�
�+47�G�!�qG.�g-D����6V1_y��xÌG�r��L�k�2���-;�6�����YP�l��Q%��p!��TKp�h�G��@�t����\#$��U�}��%�6O�T(s�L�v~#S�*4X�����Ԉ/���WX���F>�����#\V=fZ�L,~�\�F쪭�䴯l�1���`���d�&��f��7Rfv�!)�_� ��\�I��¥�����6�v����o]�������� S��GX�� �Ԡ�6V�1�Q���Kf�m5r��U�j�ٷ���PWK��eHͽ�B:�p�ͨr�w�q��m5�}���A�J(���-���0mP�u�JA�N3BB2��7z�*I�� �Υ���{�t`D4�d���bdOp�~���IN�*�qW� j�T��ۇ�Z����Ƣ6<bk���u3�����/���&b7A�oY�U�%��#|�4�_/�����Zl�H=��%X�����[:�5�e��/u� 4zh���|#�	/��9�jW�M�&K�'���U�>��:�\��gk���5#�>�Ҷ5Ѱ�>�~���]��6|�O�g�s�	���[�2~����L(N�ώ�fK9r�I d�%�'w:�"R��4���;�d-���Zm�-v`��5p�f@f�/�a�i+Q�(�ؾ�[] �$�?N<�6ma|N�����V���+m��� �3-�Z�&�f7��~ �V_i f�\0�^��: 6N�� �h�St���L�UW�H��/��!y�w��"��U9չQ{_��߿w1�#yzڠ��U\���,����?�p�; i®�Չ�F�v�2%��,�P}�(�j܋�&����x�Y#���nH�%ָ��@�٫|oͮ�nB����M��EL��c�gg(��Q��qi�/�x�6���|<�H=;)gs��/PK�����0&U�4]��i;@ׯ�ݺ�Y<#�:���{�Ҡ>W*㾓b��Z�$櫛�[��������ێ=���r	E/���- k�������+���CR��&7-�,4Y��|�ǯ�����2�����&a��~0L(��e��*} ĔP������Gw�	@q����W��C<4��KR!(ri�-�jFŮ�7����f9��N�6� �(Fk�?Y?��� �S6�L~�c�!���D	_N=|\ϔ������@��n��N���
�X|��=L3�eY� ���ꡒdߗ΍��R���~�O���w���Q2�%���=t1����)��5�!}K��;���Ղ��+�I�f�P|�����_������3�#4���s��,��*�\E�Z�ܩZ.�U�����Pj$�m�3�],n�
��\�h���ԏ�	x�I��A�T)�A�b�	�m�F�O��(P�2D�a91�>:,�[���#@v=b�˲�!�����u-.�Ȩ���	J,~Sq)�L���@\�$��U�L�����j��X�8`��FX���@4jb������[!�IU#"��kЀT/V�����Б������4ίT݊��DZ��,Yl%�z���~�D��2�2�Hw���WE�QyJ��H\F��d]~���f����G�O���/��� '~}�;pU�_1���2x���#�������(�A�I��%s$���b
���Iғ̑����I�`R��0�q7���$�R�We����0����kt��w�\G�.@���`p�5w�:Ţe��(�ѥT���e�QV���E�ʑwu�����b����F&��݇�;��� {7E<³9A��,��`NO��0�?-qBiؘ$��
���
�`Xņ#�IAXs��qo ��q=5P�v~uz��4݉�w9�FH���Ɲk8�8K���f�6�;?������Xr�����%����.n��
��`H���l�N��ˆh��|���;�'�é�2�Vq@�}'%��n; �]��9\�� ����n�:���� a�U�{OuTH�c]����v^����T@}�����2H��M�Y
-�0g�(�$��y��;���.�?�6�z��ЃFӨ`�dݏŀ�O�ͽ3uv���c�7�T��P�f$��eZ�ߤȪx=��B;����rM�os�n=�'<J�Z)/	�G���jt��;�,Rv;PE�*���P_ș�2E�:��P�-"�;9QU�/K�Ku���K�J�������I�`�9 g|'2Df�K뚔8n��Ɓ�Gw!�~sa���<u��+��iz�kV�t##��m��~m�'�h���޾cv��-Ѻ*7���gQ,���b����<6�R�z~���%�U����	f*q�.;�U�$d�8��|��<ڵ<S���a�^`1<�l�6����pō��O�;×�4'���X(�5	&Bd�r.X��/U���V������O����q`Ͽ�}}c�M�,e��40ݿ#�
�J�l?US��P��χ*h��)j��3�i�v��$y'�Uj��.�a7�'�v�$(ɀ&tV�G�x�_:�û�G�bOzО��^��-#�x��
�^���y���ë�A�5�A;]�l!Wd�ꋹ���@W��S��ϭ��0h!U�Q����*|1=��Ւ�l�pW�ѪQ[�#�n�p��I����W~z��K�;�L���	�y+�q��/@0��p��tm���KDrAv19�v���> U��C�r��j��	i��pY����؇�W�rM[��������h�]'�mj��� ΍��WW=�hF�X�N.�f��:�D�4�ǥu1P� !�S�����E����P�J����;�5T�9�D�l/�
�Y�O�&�b���K�ɫw�?G� ���DY5��O����/� ��x�.�qAWd\f� q�#���M]�Q��t���J�kP��Qp����1�{~I)V�l��5)�ҳx��'QxM�B.��;6�I�2��!����ḗo?}�b�D�l��{�������T�Ա��~����N�G�'˫�i�DwIT���� �Y����V�O���|��7$���O<*��E�e��I�{�C&Y�ӆ��YT�Y��,��2�BX�=G(�Ȃ�P�P�pc�m!AS��Fھ���;lZ�f�,$;���D�?n�#��f�R�ù�6��uF�J����6c�ok*������?r=����l��ih��4V��]эfa��Dq�A����י��/�����;V+n���Q���X����������b52kׯ���ĢG�T���*K��4�]$�#�FbI�Ԣ��Vh�,��^�&nN'��G�ޣ�N2�l�f��|�z~Z���e�`�"����f�z "��ޔ�	n8�X��C(��:�]��
s�`�i�Y&�>�G�ŝ�����Ws��%Yy���YC�R)�d���EƬ����9�tOoÕ��������w�l���� �h�[��p���)Qh�c��]Kq>@��@f��T��$*������u���6y)e��\c����U[L`J�o�ɒr�tD��K��!���
.�Ĕpeާ݊HU���A?	�Pý���e��a�=O:��=���tG97}��җ��G��|�N��Z�M�Y�e�p^�,a�#�{Ld��c��wf/_�/���bBˁ�N�n����3~Q����s���l��4�1;fD\:�-9غ���'*�6�'�8ۣ��|��G�S3��N8pF�Sv�B����G0t�I�mq�$3��	�l��ۆ4�Ԏ�=�~a����y}cй�����t.q�@&>�Ov���c��tgFG� ���iH�s�����½Hm��j���k�������ҥX����#�r��{	�0q1�i�nYsiwE����Uh�b�f7XXuH+����-P���(��.]CyU>TČ��߿:�ҽ�%H�tJ���M�ʌ��$g����Hn�+��p�꺊�Y_�+���n7#�LJ��LS����|%&IG�2����2|˃3���Awv�f���	�K��0C,������[@Ka6(҄���F�I2�����}9��SxΎq�����*�p�'�R:��(G�}�{�8/�9ׅb���2fEGl�C�V@9�%��W��Ζ����ʼ/E�6�\/a4V����DH��)����8>�h����1%Rԏ=����>a��Ȯ����K��<u�R�L)��u
1�
�C2�䫯f��"��@������n|6�[���"74�6�V�;�!� ���x�X�&)6�I��B��9��hA\X�F�%��ْD8/�lR�6�i����	���Kϗ�6	A�˨��ph�/j�����o[WvFK��>^ծ�GvY�,�U<��?�-*������;�X�-�֌^�U٤ѳ��8�b�CK���bA��*���Ϛ�UW�A6ŭ�Z"��r���r�I��u;�;�0��ދU�A�~�\	�c΁�Rs+(��h��p)�^O��
���'}>��.ld2�����2	 ���wh�֑��Cl'�{����y���-�/s峾w��4f������ؓ�M'�8�0��Rm��q��z�r�C�&?������M3.��T�'���81c���P�uA.�'�g�������"�hg[�/]�_��)t��*�?LSI�g���d{��ͯI�W�=��,������N������J.�-�i �~�dVJ=ՙl�=�
q3Z�|�{Z3��,9Ŋ�;���7K��w!3v?��b%Ns�5!-7p`��7��pQ?H�~��?���2��\{�˼%h��e�ñN>c�:�VϟV3��A�o��[Q� ��NÃ� �	�B���`U<�'��E�y���8����U=����
�+ I��/B6���� "3����6� �{��O�x��Z�8}�)�[O@����X�����	p0X~��y:�H��	-�L,��c���NF�B�v�\�����K-,:�?�.C�+[R���t�Z2_lD34�#�ة�[��؏*����겛��!�=��'��j�u�2�\`���ERx�Vn�����'A��ɩo�U�~�D[sמq��FO�����+jH����xk�N��gP�:#�m8܆���D2��͠hT�eB{nB����4(�I�'�pW�n[R��j��tt4P(�����ͨkj`&5}�Fa��s]�5Y�f�s��lq:� �S9�2B�V�r�8P�T��\XJ2��d(Pe��3� 2��$J�bF�{u����Y(En/�Vӈ�3b6�z<�_r����)��T�r�쒕�C'�'�P8���9z[7�%;�ܙ}51��o��\C�������=�c���|�s����J�^��I���Jd��N�Y��2Ue�a�38�\]˛�ԡ�Z�+�d:�˩�!�&8�f8+���⌄�{v�0��F�2�9�>�j!p��7E'.	�,7-����5Z��'aO�W�-���E(q��� ����<q�/����:yO�#d^b�>E�'���dl�EN�Vxh�4�GZ�\@�MQ�L���|���9>A��E��EK�t������75�<���H,ڐ���}'3V3N!v^N���q�5!����_���܂��WF/}R�B�b2�"�y>�w�����x��1����$7O���Oh���R������Q��H���,<�6�����mx3.��ߩ��ZD�w4Z��H/�����^v��c�go����Ԍ�9w�&���x��Kaa�2,�Cu@^�w�5$����W����2��[
��6�?���9T (.��ν͖ޏ�P ����i"�V7�E��]�핍VX�j����ԑ>\��6�,�5~HsM�����z�=����(���	�ŚoI��$��m��ײ�"=�"�&xBolY��L��`k�7nD��v�^�aPRA(7]��D�E�N�ُ@�V�aR��Kl��-R�>�zέ��_-����,{fE�u�Bx���y'�|L�S`���9�<ۭ<!�<f�b���0���r�K�p2\\őAׄ�A��](/
�،���]\�}!:�x��"^�C�*�C��!���e�Ɂ���[�C��wN��	*�Z^YP�s����} z��,EP�{�Nh#0���s��{�@�;>�`mHM�{��Ē��6�>>O���q>�Ȯ�Z���c���Q�!&<B	����;��ം�kI�����Ӗi�K���	:Ԝ�;v�a඀��k��
1����J�N��6<��&k���������Az�&@!i.56�*��l(sbz�k=˞�R�B �z|1̖�=w�g�fE��N�[�HF5�Jo~�o��n����BZ��mؙm��Js8|0*G��E<�nT�ڝ��V\��G�_&1����&Y��&?�l����A�YT�z�Uދ�ͫ��r��%��l[���]�f\���땭.�ؼ�)��;DJ����P��n�4�ˌ�lO��5���/�_pa0���0Q�Q�SΛl�a���Zt�~T���F��dm��������)��r�|̰��A���J��,sύ�O�F�T�k�jg�$�}�n��� ���o�s�Ȭ����o�z�$��"%M�&�ORMLC5����>���� &���F.�
���V�+7S!�D3+I���W"����,P�C������ôf�'z?����d���c�P ~���\���,�Cdq��������8��&pVV�j�
#�� �LiP�z4%��0��g�C[?q�����Eu�͛���^��aG�]_��$ɔ�Q����y��{���ߦ�f,}��w�YBm`����+���#?��uO﴿[+)w��Z1�>o�6=@��Ǘ�ç�1.���u1\=��\[�<��s���gˋ���/M��2���ʲ�?�~<R�\Oښ��#x�<`1l֋��8О�&&�	삽U�� Zw^�Ā�=�E�����P4k&�SK�ٗX��h7l�ُ�91_��Jz.��e���8�'��-a�#5H���O�b�9iǶ#S�in�/ �4��t��خg��ؖ`3�X(��o"!��fL_ ��gaF'([�3��?���3���zEV5QOG:��{��_J�s�BRQr���3Щt/�y��-t��o=�R+�#�[P������b��R,��������#6T��4��n��@V��3>�����iܯ%�|ɑ�U�n^bw��,�ƐN[���mM�)w��0�xRX�ݭ�j�ƔW��D�
��5�&#�a68��a(=���wj�)�:�G�CS�/	��xfܓ�-�Z����W5R{S�}L�5)���q���*C2� ��S(d���N����_�[�$����n���.)e�v��IQ�MKv���A}�b�B�`E A�K�p=���]�Өi�E����N1qt�1�4�X渐-�iEN���$��jV!��������\۽)�A�����\]�/��ْ����}�wb�)�A�#�w���J7�&���M�D�`d��
8&��:�o���./�r� ��uR+rB��I��܈=9���E�»���y��Ռ</$��[T[��(�*C�Ih�cL���7�[�ck���nq��O��L�i�b���7�Ty���Ys׮]���b�BND���U5+3�����Ann�]N��_�5!�9�t���yy����Q6"���?�Y�"o�/�+���>�P,�`G���`&��z��?�K�v��ˑ����{��/�����V��b�l�����Js�eM�2������M�Ur�%~,yaZZ��K�]�=��(4�BhhXY ��ȸ�ɛ����k<�sx%1��Z3IȤ�U9U��7r�=�ڤ����~��}z�������k�HZx��jB��C��V��z�����i5��/��RN�`[R��u!���(M.��ޑ/�p@�@V����HR��1���7I)?��}��pQ� ]�xe}Ρ,�oͳ�	f�����_�S��Q��h�P�c�x�*��9��� ���49
���	2������F~�nQ�a��"�Y�_�l ��#PW�Zz��rJ�aC܌X�B�K��ZcE�m�8���P'��1��oixY���E�jC��ou6֗Fi0��ʨ���Ve��9t��D��'�:�~��E\��5�F��/
�����'�� b@4%E��ā�W5ۜJX��
��	9���h�1O{���Gd	�Xt�v2�Ϲv�����ͼ��V�SG�q�;�R����=45'A2����%܏��^��4���%��t�=w�
g��t��wOc�̤��5b�1�&T�j�o�JU�*��혔�+�t.j��(��/�8݁��ȍ*P��Ӡ
 �(�Y�{������4��V�BFq�����!�
ρ�8��f_�Ϊ01�&p��vX?���Ha�ß�\h�~��[}��7@2I`��j}2/ D��_���#!݂ V$�8�U`���`�]_� ���M�\�$:{���h�\�DF%S_ꙸ�S�O��V���F���)6��0��T(�j,�2>��ɣPm��T��JU't���8��"$�x�U`�Y�(hͼ	��D�����Lƿ�oA�eO�z�|���$@}l�X�����M9���D��pJZET�x�tI�����Q�n�D����R���J�Q�c��=g*թw��b��,�Z%�	,�2��2�J� �g�نK��5{iK�HP��:��4^"�����_)�_�g�8p�9̀�g/�_;��� V�!M����>s9�¬AO�l����^���G'��C�O��p�jp�LY�^�a�!ًAe`��"N�q����zaa�l�>�퀑�m��,��r�j��F���z��Ʃ�{AXC���ל�!�]:���S����;��˥}��T�d��E�z.S6��SWGDC.��:rY
50(<�HH_��2b�B��#!�{�z���q=-!�q�6��V��B��N ��(&�M�ǳ+�%�t��*��1��|'�%]��6��hZ �r��rP&%��2^�`_�z ���
��1D|܂B���5K�/�;����(��D�*rki8�g+���pr��]��"+5�|O?�Su���y�gL�^3���.6�E�drm X� �6�_$�dV�WSJ�����9
��D��PT˲��[�q��5�';d�6$�0�F�h�G�ŗ��U�Io+�U>h~����������D�:���x���ίs��)�<	/� �Ǻ�趸�
�<��h�/u�Q_<�����+���a�����f�qŊbC��U�B!�M��n�n��N�U-x�W�ގۛY�ܠ���[�8���A��y��*KY��Ѭ�w��,�������?�<KIf�����$���D�M$!��I��jZ��9	e �ھx� �ζ���J��c'w_�N�_˥��w.���}b�Vn��. �H�Ҧ�l��\�#�qG
�������v?u��<YP���l	� k�FD�i�R}vT�-��,2��mf��0�?�P�ғS�����\�{i�k��"Bcj\��^(�V�]�|O�����+E�N�~��X��*Y}����e;c�?`h/�b16���FF|�5�H<�y���T�Nz�w��Ϫ��v����Gⓛ/b�}�gE�;9�,`����(*�[=���������79VT3�9(B7,��>�kt���s�]UɽΟ�xb�t��M/ 7sc�P�&0�8� ��n)Vu��y �)M&�l)��VRgS{_'�Q��_=GIi5������&$���1$u$
;4j/B������ P�:� ��I��߲�A��Q+r��,GD~��㛽cQ.w�9�4�|R���v()���%3;�3 �b�����w��#���3��7xFb�����gH{�W�j4<���rґW:���Z���!�/|�Ϯ���#A�'֦:@�3`�U;M9��7Fe�Xz�M���ڵ%22o���&LU3���]_g�=@��B��BX�4��7�]Wb�cZ=�$"���=�8�`��������wS��\����"~�)�b^ID�z�k2��r�΃E!�3���y]�.~�~%�`+�d��f���������)�:m��'Bmp���iqFע�!��k����9�E��wQES���?t��Uʪ@�@�,	��~ �x��K����a4ի+�I�8�|�S I�
�E���KoLzaB���턗����ݢ�h~�Kms�^(��) ��77>K=>���¬'��h+��X����v��'J��^sN�~�/��+t�#xx�T�!O�E*�a΂iP�H������!,�^刢��QwC�):�*��k��]�/��K�	(⠁Ȏ�\���%�F��~W��^��]Y��J�!C�Dy�rtv��G��$�}D�m}d'�;YlDqwcaC��QI?,��!�6dw<���n��زŬ��6xY��!_�
����v�C^�'/QX
��ɪ��+/̶��j~�n�<(v^��.��}��Nua�Gg۟W�g�chު�DU$�Fv�e�D�n�}�^	�������<b9�5�=s�'�0�ԇv�����L��k�]'�C���.�嘡_,�a� gR;ЮHI�t�mU@`y��-[��%Ҕ)��>QRFo!K��J������j\�����A�ň�s_�[�W��D��j�o4��rbA��!d��:*�=���uj�z���O����b�H�v�}��I$N�3�:���o�;��䭃��)�:��C����o_Ɔ����1�Q�Y�1q�L���4=��j��G��Y�09؀�����s�cEf���}RQ��V���Mme����\���g�0Lm���%4�D��w�#ʺo�*m��0���I�XQ6!� SJ@�p��OG���-�.?P���� x���:��<[�1
�]�!�ԏ=�[jl�R�MH��7�1�+	�:�}}��� ��=�AM�]�J2�+��* NG�Z���)�����Sm!�m0c�3u�ME,�E�J}�]���M���� c�C����UKd����\.�K��""l0ܦ[('E���!Fd�7�v�]�32e���G�nMT^8�#8�{�e�XLR\�3:��j.�<��������o����EJ�
�'ϩ�w4���%k>�P&A�\�>o\ϙsQ�Vo�����I��
��w}��L��Y��?d��:t�m:����L4m��:n��C�hB������h>*8l�U�4<�=�)A�H��iVx8�O;�TGS-�*�]���]��.����đ>�q$Qe���*�e ��?I�
?�/Mh-���V����6*o)d��t;�"����}*���*��=�5�R�#cV�z�)ـCH�R������w�L_=׌�zV�Ȯ��]����wB��tW�E�[¨�#����p<ݬ*�|B�7c�v�}g1�P.bŠ`M&&iJ�.	6N����X�t�m���q�y�d�O|�z*J�Y,�D$R�6��!�^�-���,�(y�|������?B }
��V�� ������l�1 �V�$�U�یO�A�'#���<en�js'G#޷�hW3߭,���A�n5��nwQ����)dLӲS�*�2gX͵�\ ��}l	~�o�A&�1���Y�����U3<�B��u@�Z�S	�c�m�>���&!S��#H��S��I5��`�5��Eh�0���3G�����gYW�|��z���C�e�ܞ4d�fׄ�΀�U=4�n���{#}�yNy7�^��j�O/��_��$͸�-�ı�-1t�#��䙹�wagN��~@8T�z�qrUTg��8P%ˬhv��������s&T���eF�gd>i����ۨ�ڤ�^�¦qڀHQ�l�,af�W��Y�_��i���m
�:�N���]7�^�OeS-�@С��E�!�< Hq�B��0q�/<���ˁp�W=�-MJ���(��R�?��.�7�,x����[ÆN���2 _�Ê�X� nV��f�P��,q�n��$Ct�����Xz�vZ]sLX��N�2��d4Nj2�Y�0�Y���0��U�ק������A�O �nHx[oo�S�M�WRI��e� �7s>��H~>maM#5}>r�K(`�r{��Mw���ХH|�#g�v�D�y���nXP������yTu��d	�.io(�1�6L\ql�D (h�i�ʰ�Ey�]ˁ�܄�Fp6{���we���D�I԰�4�������^)�5�-�x���]v���\�'��������Ԅ���2J[M�6�������x��-��Ղ�\;l�+�+ݺ�89g�ϲ�W��JR�\��½Y��i�_���6hF��6>wkC���ζ}u��ʙ���]�e����{D5[IV0+î($�7���|)>$I>����n�Y/6��S���;E���Kl��ek_�PB2X���+W�|�t��[h������zJ{(��V���|Af	��8�֐3<�F�<܄�!��4$8Y`��"��Qiڬ�]|��/����d����@�o�#}`���X⢲�.TBMՠڇ�cП�`� ��; ^&�P y,겞����h�ό�z�+���Oh��w�4����{�ʌ�p$%�Y=[����)�1���o�~�{����������_Dn����V��B� 9e<�j����u~� ��]b11a$+|AP�}SL��=jQ�7�H	�9���*	�^9�ʈD��?V�<s�{�w�.&��ǫ+�zD����ʲvzqn����n���2�9�b�n>dt���Ox^�@:T�̚v���;� 0�X��E�R{5ձ��`��{�پ�;�0�Jro���Q��"�mʜwu�	�`�įQ1Y̱�����D����M<_���w����/q�b�#�]���2��YNGZ�����n���T����γ� w������8�>G���6��(�J��c�M�hK�i�aD;�K�d�B^�Y<i{k��z�	���'֐�7��`��U�e���&SmQ	&_ I_�5W��4
��օg����9��ْW��#s-�����-�o��ƹ�Ȓ&�r��o��~�X��Fn;r�x"���5�a����Sɻ.�T>'�F�iTs�Nec}0���-mc�[�8��Jg��.��F�~%�j���u��$'MOV�dF�)�UD��}iB�_�nB���	�w#�͞��9�Վ��m�Q��W8�^maP➻��F��b�<|;@W��%�+��p��� FX�e�K��X��M=��l^bb��y[m����0I��=s�X䚳�{Y��!|�e�=�)�eH}�c�K�������7?� ���9��i�L0��5;b�d�@4��jQ3o(��Q�������̲�)&yt[~5�k��8Ⱦ�=�ۺ�@F"�6���o��l�z���x���'Ym�83X�ϱX>�=�^�A�1�U`���;�S��Ē]�L��Jl$��o�!.\X�)�ʋ��q*���Ϸ�w�\��C��D+��*h)�Qh)�W�Xs���Mn�T��oBtn���n��â��I�^������[�|' �Ժ��Z�c� G�?%�N��#���sEѷ�&�ώ=�@#��铬\.� ��
��t-Ȣ�=�8��,ӡ�NQ��N��|���Lj�g�� 9�Ƕ�AMpްj�O��a�&�ء�����=�G����*����h�G��Ün��BkDQ��F��5��+�|ݗmV��es��E�%:���s=�ײ�2
�s8^��~l[�y�2�pd�nPlՇ10;�K��K D�;޺<����,�xD؜��7E���MC����&jԚ+c���z} �=��@��I��9{��$�S��Do'��h���g�����{�ؤ�&�Joƚ�Ӑ�1\�7�`U�rZ���(9a����F_5;�@�5Ŗ��L��o�+��9{��%�%TS�����o��ʰ��rX ���7�-��?i޼���'�����;���R\h	�1Dx���Za%PV���o��uG�i��#��|�4)(?��2��ϨT���\|_�H+\�g=��RJ�B�z���}�}W^N��{A�]βk� ��]&��[�_ �O}��*?qdr&�����aJE��N�h���7Bm�޸�T�f� e���z�ߙ��$�P{f|�3�Ƒ펨�`�#���)E��"zBw�8�*�]� �yJB��&�dQ(b���C��Sv40��͢��A@aF^k��*�J�]��qpm09wE��R�+Ȋ��k,L'2� x֎�l��Z�)�^*���4�4~���h���G��>F��bx?�I�zhfB+��+�9���N%�D�ep<�Sg	z����OO�Φ�sO/@��wL*a�sA,�V�v˺B�{��cr���Dl�cջhM	Ᾰ��1{��Uǫ�#q�-\i�T,��)`��g�Y}��2㥝��̊y|�P���.�;����'�y�v�n)
��?�@H
;�Hp�ڲ]W���7�V~�;�X�������*�j�!=hO��[*"�w�b'��vٟa�`D��¹O����� ��R}ϟ�n󴕂���
���fu;�������m���]�dn|�(�8�7ְ�u�N��~|0G~�?�w
��#"d���*���oJYk�G{PE?��r���	�mYT&(�8I\Mn�?�R�h~��� �.�8C�=��',���V�R"&��y�/��Zk�S���zGx'�����`�G\N	�n�Z!��yA�!E%'���#1�r�yi���]��M�Aw�h扖����̋˾��_H�)�ǯ	w�|� r8�ͳ-b�"5^7U�,������s�z��<a�B���ȥ0�C�aE�����ǹZ��G4��8�R�F��-�b�#�</1���S�A3c+{nv;�9T~g��*錈́��!��Ћ�m�d�Q�!�����g�ZAEV�{h�����>	�LS�l�Qe��7H�	"2��q�c�&��Cu�������%�P|�޾ь���o��C�^���x�mr.�BwɄ����č�k���T�)��e�v6�q~�G�H�d&z7ݩ�S��{xo{��Ώ�f�	_R-�_W�I�
AW�	�����'R����gd��	X�ي�U��(�>�C�%�-�;��#�����1�1�X��I7���Ӵ�,�B��!�b��qD�+����,����j9Y�	�H4p�X�D�����ߊG�ǽ})��k�_L���XJ	ȉC[�AlYD�N�?�K*�`;?<�c�2G�:��ƿ��k���B��`wćFc�53I�Կ����ɫS�#��Ք&�[3�F���X�>�@C�k���Y����0��=S�KP4nS�{�J��M�2e�)C��f��c X���3�?�"Uo��]`�wҜ��0������M�8ORP�p|޲���M�<��&'| ^`V:����P�Y7j� 3�4]/-ك�o��?��Ncu��7'|y��p��l��b��0~zi56E1.xU5���t���u	x�?���9\T[��%])�>�W�qԄ������i���\�|��Pw(Ǻ���HF3�����;p|*����t��\AŦ�0�]����[�[����8����*g/�$!�n��ϓ��o��G#�=ko�U0����F�oF��.�,u�
��-A�;�%��>ӿ M\�V�&;�����z�$*>p}(gF�X�z�鄅Z����b��lRlu��o�q s�w[U�i����{L�T[ҹ�`��;	��7�Q���f?�' 8�<�㟽�81&s�
�%f������k��׼p�b�p��N_6�
�����鲟��?����;�ND��D~ahs8!�3�^I�_6Ӕ��kn��Sʑ%���y��IǼ�5�عZă����s=j�+�0s�����b��]Q-캃�I��`���$��e�����E^��3z3H�E���p��<��8̴�߹���������$e&�L\��������5��lL�%M�6ѵ����/�(��\��b�C�wb�&�㗈��CT�6�4B%�ְKwe	�f�T&�@��l[-�R%�ZFi!p��T�c�����E'=���5�Ց�~]���e�>��Ƣ��R�+�O8��(Z7;f"��,�F?#s]n�%��Y�"v�m�RsBJ
�;��8��	|�:x���L:
Eu��_�V��{oð�H�#-�b���+g
�7�U�>�E�<���$󳢄Q�(�����L��$'�|�}��P�f��M�~;ǿ&��y[GY�}Z6�`
��?�{���� Ry��ޫBa��,�)I��|�O<�t4\y&3��b�(�dR��'"���c����s��0�7�Ǹ�A�&c�6�f_�bȽ�.
b)�7���j���<1]!���!���n�_��B��5��K��w�t����5�:�\^�!k.E+u��X����Ն$�w�Ӫ��f��v?%o���(������c��� ;h�W�ȿ�Q?B�.�Y����<��n����>O4����M�^0���c�=�X��@bטr�R얅tJs+[�n��2\�����<��oess����QYqB	n/�@��	Oc���?û 9?y���u�Rֹ)�`��eγ��8�J�Aky�AO���*�W��]P/��U��݆ܾ�5�������@�\�:(����I��k��R�����/!�w�&-P�Sh�1��]��A#U��"I��Kln��~��q�r���i b����h>�#��qM+5׹P$��y@��������ｲw�U���QD��*Z����"B�W�&��VpIVVS/謥�ƃ�S��nfV7t7��u�g�MݨF���&$1.��r^��:���1���#��G��)�{�Y,���?<fݔ��^}�i�0m�i�Gx�##�%$��ML���u��2����$���� &~oڞPҴ3kF��#Ļ@j5m�9Fe�L}(,���G��'��/nT̎v��h\=Vۇ���O�tOR�pp�I�T(����i��]^����iު���t��sc�BA� :��VF��q�P�	3֯����~/ߥ��*��g���X�1� ��D��_�H���8�汦n2�T�}�4C��}���d�z�k(��'��c��xf�A�<N����:�r2�!��R���jIs�3�B��2
ЯN|%��� T�hG��߼�:���Ł�l��np� ���4�(���&,�s���Έ���w'��8�ʑj�.�W�4|uV4Q��uZj��V����l����{x�)g��
��|n���*Ed�LyT�h@�2���`�_��@@na�5����3S����:]\��q����s��&4n���΄�"MMJ����m���2	����Wf�R(ːNJ,
�1(���b%O₭P�.,8H�?�3����$*�6$�p��޳�<�4���N�9����໌>_���߸�]v�E1}8(��zN�r6^�mk!i]����Űy�]�jb�f���\��%B�JL~w�?q���"���R۫͜L�]��6��R�sؗR޶�I#���6}f38��y�b��v��v�z��4��ϏHW|�Y��{��,�6y>/V�^��n��݃���q7���kEeԙڐ��֝��M2����D��Q.b��^�!�-��	1�E���)%92�;@,��(8̀u|�_]v��f2CMx�l)׻�̬I�5�
�8��,a�5�B�@v�?�d+Qxա;Gy���.EBdkh{�MjG3�pA~Ϋ�g�o�ڞ����H 1r��F�6,k[�b{���ދz\n,�Q׆AчY�6{^�uYLm���W�2ӏӻ�6�-4NZUm�0�6_��1�r�Cs�|�9KČ����/�����K��-{�����^|�����"�b����2��e�jkLN���9,!��h�.��_�����sf�cm�+��DZ`��hit�A�r�u�"*b�8u ����1t��~oPlA¾�4�1'6�Ou�;G�F�0֜�/'Zw��Hŉs��Q��L������o��� ��װgL�.���2�}6���i��Y}YM����}�	��|4]#F�S�/�Dt�+?��-�J�D:�RF4P�}vu_��Z�v3�3��+yO�m�I����RN`�Vk5���HKwh�A�Dλh�[��Ie��5���c�V���iW&���y�.E�
��|;�
��`R�$�)��ɿ���W�Ĵi8VEr!D�����O��?M���Z{>)��Ӱ��pf%<LV�2s`���݇���m�U����N/��`��ˤ�-�����Bb$D$[����s���q.�:�E����A�i3Ac��[q��`��5��-e�_����c��٬0J1�L致q�̘C���C8��,y�$s��q�_y�b��'�Ƥ�"1�U=G�;}]���D���ܒ?X�����~Q���ڔ��$��!��ɳ�|� :�kw��?Xy�`T� ��"�j�m �GJ�F/.�To�����5@��gF��/�*X�:�2ɇ0��𥮱˄�
ᦶ���C?`τ%� �Y�lO�T<|�Y�+G�݃���x^E�_^��sQ|�d�TCV��wz��_-�/r�I�̩I�����j�!��F[�	�o�fװo6����u�9ף�%?7a��Ev(ܬ���ݸ�V#��g��vz"��p�E�������aM�����_[e�U�!�6��BPO��8��xH�����7�L�>�z��z�#�I�>Ҋ�y)j�~��]/\���%�`]ձ$&��;x����6E&�a�D�$�!�����X�aSY�u���	>�t��0h�mW��&4EMg��F�X�Z�)0�h[ L�0��|��5jxS⑴D�w�  �`�V��2�8��V��A��ѷ�b���M�K}tp)RG�j ]�҄�N&�xq�Ȉf��l�AC��G���hj��!� �݆�R�j�2���%54e��������L
{���t	ݨ3suPH`�]uH���ѐ��?�s=��2.p���8`���"D�T������L���g-���/ `�[y�zub`Ȟ9�r'4�>�÷6:�Z�	�_�Rsl�rۗJ�KJ�w�G�=��v������Ԫ�J�f�/��V�3����,��-@�Y]����<�y
�`��d>L�M����̸K�Û�h� �����9򕷢����d
�7(z���o���c?G7�}�3�h�I�Ϛv�Zu��3m���V?z\�@{�k�0n��_��h�7+�&�6_�zۈ�R�{L�� ��w;o���e���7궬ˆ �p���d�K��-n� ޚ=��W�B��Ճ"�k���y8�]��F�+n���3�#�کv�a� p֣��[|�M(��Clu�"j��A��]P����xݣT^��J"jT�K��9��x.n(��㚃�_v�xԛ�d��bZ�j�4`�֮���q�D)��� @4��3;%A��?D�� @T�7P�6v�#:@�|b0��?��H�(�AU�E�� ��o��b��|��qj>O�A�
t�_Y�q��}"��:Aӻ�@M]��ToX=��s0��J���4����/�����M��l>�p��&�[y[�f"�����g0|M��{�T���5=���9��k��S�_o�z��Ɔ��4qh��c�wvr�׻���F�Đ�*uֶ���_�R����(_R�r���N�I2Sk9�Cu�8\����CQ sS�BC]���(���QHy�qL���Qk����Af��!Y
X4�������	(|ؗ��M�+�:5�f��B���k����!�(�t�t��/��n��:V��UPw?XM��� c� �v�^����@��Z��1�nf!�UΠ9eƉ!�J,� ��Ɇ�g��i��h��U�푀]��[
1��H��cq�}4n�Oͺ��0�w7	��]u��c0ե���}r�fcH��4�ma�g�h�[u�-���2��qxf������'.�Pt��[)��m���u���->��0F;���©�۹��&�x��4�z�粁�X�	��5U�3P���U	þ�
D�������><1pwϐ�)�&��/� ��yL�r��:�wU��a�,.�d�1�K�S���/G�N��P�Q�!h!�j��i'��RIs�b!�$l��)�wɮ�J3��坩�_bרۢ��Æ�Ղ�L��y� ��W�P��Y�T0p���}������t%�6f��N����&Ay�Z���	����2"³@`�jt�؝�*��t9m�x2�ۅ���7���t����.��C� �L�:Ku]i�ƻqH��RĞ��m�SϢNe
N���sx����t��e�����%��>�|�}���G	=�3��� *Rs.(��\b�[���s.����'�X��r^����k�-k��*]@Lnx\Ƥ�"[��T��{��@��Nm�/M;��M}��jM�ﾳq�n�y	2"F�F�d����dP�x� {L�b��w���Սws�!T��h����0�9m��n5���l�ﹴ�9��c�޴��dKa8nE���A A�H ����x�g�j?eD*5�,Ԉ��zᏘ[j�ٙd�
��,biL
�_����!��X_s�7���K�8�7�&�цd�e����f���KM��AW���Z��tl?2�6�R�뷃�T^-1r`7��`\���:��P������K�u��`�e?�2�]BӋ����������Wߝ׌4C��4�H)�9�i������H??����ѓW���o� �������W���`�U�F���I��:����{��T���4�9����A��Y*\�
A{i��u��3M��wB��K�8�ǐ{���G�f�6d$�����Τ@v4"�AY訙L��Df�"��6:�Կ���J䙧��c���x�"}.���4|(˭Z�� �f�3�۽Q�֢�P�lZ6Kvo��+���Mt�.�jq��Ww�M>m1�N�G�s�?L�SZ;���$x�i�O����!�x���CR� <�'L���07;�w!�	���(\���pZx�E5��B���ɑ�g�@�,��p��~$�DJ�Z�E>�?h`�y5#�#-��1X��viF�D�(a�I��F��]N$
�	(
� �=&U��L�|"1�E��ԛ@w�����q�L58����5�����&�61���3�Hl_�~�����1�i�=Ј`[ٜ�k �U�h�yν���0�$X����Y�]��v��x��EeG�A�k�[��4s���:꼠k �;�$�ښ峁j|㑪�jh��uh��}CV���T6��ϲ-�K��!����_Y]�g��O���ed�$�I���B�Ii��;��@�e찶��MOk{��`��C�~M�;/ut����ul�D���x��Э�`Qo�d���uQh¨#�4+w]ѳ�#�6�z�/ �v�HJ�,�YpTg9�h�4���O�������#x��9���Wǽ�v�8������+Sx+�{�R��8
Qr7��;�:��q�K�+>W�ٯ���V�	�~B�<x�Z��ݞ�/�	�^�%J0���Xm5K?�¾��l�U���H�B�2_�
:���e�����#$�tp��*�Bc�=��B�L��Vڪ|�K���q\�"E�FJ��pdrH�u����ͱ�S��=f��}�^��9����2F��7A��y��7�|d���E��)����f)ͥ�Ɯ;�b��o�}�S����5w�~w�>�#X�Ԇѥ�G}�ri$�U�Ʃ���[/^� xm�5cX�q`$~�%����+�p���dh��ȴ}pN�ǹ�@�[��{U���fU��FÐqy��V��g�ԢZb�YU���<6nӋ�!�o)F�Sxkl$7H2
�	aM=�˾�m�c���>���#	�kqxb��z-V���p���Z��x4��½d��j�'?;���0Z�U�T���P/���5#E�T	:�X��� ��L��O�d6������-�yЀ��{u��!5��a��yG8�0a�a.�YZldU�7�1�ڏ�=��
��s��Ƅ��bݢ}%ׂ�i��f�ܨ5���&�WQ<�2Pl�RC�����`��$�5س� }�h���u��NjZ�LJ($=x�)�B�ӄn/�o�'�$�ZP��z��Z�RfWjXw=Z"�O�$E�|�^_�b�8�q�-(�.�hsU�Zi�{���i`L�� ~d&�%_G�kg qF�ht�]ך�)M ϵ��� ���#��%�������9�����$	 K�+��M�,�(	*���2?i.hV»Y១E���7l4b ��uv �l�~�I ߯=-v�l�¡�����s{��AƖ]��Q�b-f��K*;W� 5�[�Rf�5�w�O<�n����B:�kYXU�إs{/�'.���DE���}�]��t�!78��zJ||�A�$�//�h�A�Hm>{޳�D���[�>���ݼUd��q�-�y��:8'ߣN�%E�� ���`f�^}|�
6TP��]69�4M\$fa�&�t7����Y�z��?�i����E-�éV!�B�M�
'�Fk]�*�{�>m�?n���~��T���w��:�VY����<�ڇ�.n>����g��>���db:��pj�Q�G��X�<��<�k�@��Ӡ�)���4����y��戯)kY=�LLΥ�y���w�q~��P�6l�6 *�F	b���;����-'5���]�F~yx�\���A�dO?���ح�ʸ�h��Q�@���w�Yb��S�e�S�T�ZR���=s�~a* �{���8S�{��a��ef�Xڧ��Ɗ�l���e )}��mWMv;�nM(K����<w��-�eeG��N�m�`x���)"��o��`����7���TV��A�@�c`�/6�D(�$QV��,>-���⑱�fU�����ݏ*�'~h>n���.`�u�-�/yf�5F�]�P�2K4U~�!�d?
P$��g@+d�{�{�MK�x�Y�p����5��������Ib��8� ���D��%�[A�ٴt���������6�����h���\]Z̆�W(F #=�Hj>�Mӗ^�����+OB�2�.� �;z�I����>U��8�:����Ž|�2I�B�x���o�Kȩ�-e�F1O� nnZ8V*���*ʔ_�`�"���3��%��Ќ����-y�m2K+ޮ�V�:���l��s��*}r��,K�7c���]Ń�F;w��#��Z\.˾�C�H�w��>N\D��~���yğ�5�i�m�V����� ��_z�u$�BoG	�.i	T%��	�J�\l����4��>��H��.w���#��Q�W�/C�-R��6��h�{t7�JAg��/67��=�F6��DKހ�6�tq�{�e� K6��?t���Wo�`��ӛ�A�77�k����$u�.8 rVӥ���Rm24����Ɛ�e�����d߼��Ø6)��[#EB_��I�ը� BP@�_�0VM��P:Zm��Q�g�1�?8�W�X<A�|J�uDv�`���V�f>�s����人_{�0�j�'��17d'����P��Lu-h���9�t�HyC�!��%�y��aT�O[�k���YTկ2���l�	���E�U^�>�R�=��u���W����3i#����)�mY\V��RB[��J.�3�=%$��n���S����H�w#��I\���OR�i�C�w�-��QTr5䶲L���mE7��ɓO(��x{���t#șXtH��Q�J�g�͖�S�د��d�i�*vٵ�.cX�Zx ~晣������k�}�W��s=ox�m��D/�� Zs`��ft6I�I\D�t�k�]i9;�($���%���+����J���.�ḓ}��Z7��+2jp\�`Ȯe��bdn;D=�4�&�(R��{��F+�^�J������9$KZy�l=������mj����q�T�V��\�+Z�O,�4JUQ��k��l�y>I�� �O}�xWn��]˩�Q�x��`+�	���
�-L�Y��M���BB��Fx���3A�9tCy����Ve�;����M�ZdRv[V30|+�\�/���\ȭB4�A�v��S�)gD=@0P����׵e�I�%~�\�V巚8�0�y.�'-B,bʂ�,������s�@���J�e�;�I��C�.���L��2jÂ���������I1cԇ�N4i���\�~'�>7+k�8V��߈ߣ"���s�?�?��ч���n|�l^n�_K���,_�H�����?����"��>҄��[�HH�����LC#��n�
��nefn��]D�T~9Z�`���X%|~��$ӆ�\��ъ!{c�N�����N�;A�} � ��x(�E�%ح=��87��l��s�����f)L���)ɋ��i���*(�)�.+�[\�L������U�`I9z�^_?�����O�>�J2�7���� ���.�R8m5��~�nn$#��bU���);*�	G�]�C�B�ް[=�4������ǝ�b���\V7 5�Qf��L���CC�݇b���E��O������OPTղ�
�� -�H��M=�qY�-M��<�F���`)'@&�Z�yX��JOb�'#�D�U�r�Ϫ
� 5��Z����<���0a��/wu��so�$l����U�j��~/�8��?bAl���ʹ����?�L�.�Z�=��	��+!��#�4b�D�Q�扈��^�lA58h��1x�!D���*zT<�3��Gd]��±q�k�7ʹ�e�J��=����7�>��\}Q������i ��[�e��y㻊��o5@���Y`��m��F)ɧ4�Q�O�LD�Z�jMQ��ě�dƇ��u[b
)�noΦ��.�k7k��/t!݆�u[7B��Y)�^�j��	�7߂��c&�r��r�Ӥځĵ�R8�ӆ��
T�m�Ӎ�
4�Y��i%F��%똨� ��T��5lT���	Z�Q�2w�6� +���@���<�]��~fi����58v]����q9��ׂ��\��|��P]<��C~�G�q$��8k.��X�W>�Cod��꺙a�3Ռ�@v[PxD�'��/�H�cS�/Gc?U#�b���!�%$K$��?r����'j��B���'�-,n�s�I���V��P#�Xks|��}�n��'��s��Qy��u��f��V���3��EN������;�N����8Cp�9#��D�n����W�3CJj`r�{��_�}tH ]�W~2�O���G�_�ՊO�м��[�`/J��%����$����q+R^��r�w�]��c/=�ֵ0��K�- �Ňߝ�׽�vp_���������������y1���sk]5�T9��b�W�k�r�]Dl��}�*�]���������B���-�t,��%�4b
�~�p��5]�b��`V�u�Q�v���i�xXB�P	$:�%>H6��H����^��ۛ���	�|���`_e�^4�{�2�-8m\;��,r\�ˢ�ˇJ���I3+o׶';�`�wP�U_.k,�˳#�I@�fnΙ ��_�.du�K�i��������CJ���L`�7��x����-��V+��+�G7�@���*�q�����XBv��_��x*���hJ���{'#,#�ǂ�����U�;��j����|�@U������ͳn� n���!�?	�{����FЈ�?�;�A�պ��a�<���6}R�����
>�c�5�&���7�kCA�kE0�9��Ƕ��sc.�J��P�����̭
��;m%��b|��1vmaq��������;�s��%���f<�>M�O�%�>�*��㝞�¸j�z�+#xlC��ǗZ�<MT��!����Z�H�=~��XS������������:���vIY�2!t<H5L1X�
�BN����UZr`��i�珳��N-0N֘6K��H���`��^�$m��:]�y�b�!EMļ��08�x�jFEFc��~piv8o���*n'�Dfb�*�{�
�3��w@�0H��{n�
�I�xN����-�[L�~�L<��?�{�rE�ӂ�+ �%���P�D�![qB�s����m(��_�+�T�`g��U�_]O��8x�΢�M�����sX�z�	٫�[�(�?��.�H]>oN��$��c�� 	�^���H��3h��,����4��+�1��u�l'�.K�����{�n|"A�\�=�Μ�� �a� dNs��z?`å�!`���?��:P�5R���2Kg��sm�S��}�eڭ�l�Q"�
R_w��2�4~e�����7㶤����H��|����	OJT�##�)!��B�����=C4���Ǖ�W㫾�\T6���;�!�(ܯ��P��f���'N��.�%U��G'_��9��<I����p�lDf&Łώ��o���;#��#�>f�k���3�{w���J���������	�b=$Y�(���� �nh<;�-���H�o��^UK��(����Wjp��d�wl��v�ɵx���*��:�5�����e��WǮg�$S�`疰DXU��ŀe�l�n�g(Q�4��0Pyy�2)�����n����o����04k�)*֔8d��qJ)*͖���`�ل�=�$!d5_Tݚ�')���ײ�֭�ۺLD��C�v���Y�{=��� +�^L��b>nɲ�s�����������X{��X�F]y�C��М�R�MԹ���c��Y�%#�;�Թqo�K�w��<�|rװ�D3�!�P64����~k�>��;�I}r�_��2J+��K�:��w$�(JY�b�Q�Ǿ��S�Z?{=��hvj�c�J�j0h0����G�JiĬ�[Ћ���h/�U޷��k��=.q{�TƔ�ٓ�p7=2�'��b|�����#�РD����8'?���i�;(�ow�ς=\��]�d��"����މ�VVj6�_��|���qՋ�iʈq��;�W��)��?�iί0M���KA٨,+�&BH����;�a�������)kn�uq�p��af�)��H�aO8��Ls$G	�J���&�%�/E�D���Lwɾ>��JR} 6j�;?��$��H'��w,&�x>n|�U������,\l�`8|�d���U���,�ǒ����H��Vw�=����O�V ��4��^�*���v��@�S�(�1=E�%&R��7�K�0��)����+.�&u�_�:G�D;�5��c��QY"Z,t)�Ac2�]F�*R
P�� O$�X�e�x��6ou�j�Ov�OJ1��!t��`��������o\c�6Ao0%����|�G�[����.ϐBi&1���7�m�WLg�{����x�/���ژ�7�L��h���$���꺺AF ;�۽��������XD�)��y�q`��qw#ŕ-)33;� �Yb����a��Uq�8m�ai�,�RH�<k�ˀ8x:{�ܫ*��\�o+(>��gn��� {O�=*$_NgD��/��Ї�]�Np&p����d�E��9�џMs����/��P�mK�D��C����h�6���������䯄h[KG�~��ۂ�_b�f��O���,��(nC���/,�95]�'G��Z�����~�aU�S+1Y�R��w�L��8����d���jd���*�-�Y�ы��P�]��#��[B���VՅN�����-R!.��vQK���-J	�gͥ
Ń"l����6�8�%��\�g�u d�b3��'-2�O���Փ������W��us�.���Vf��N_�p�_k��W䳓a�՜1I�ߤ�!%�\�ŏ�h�rN1L����E����G�u�'�3�B�	7`]��N9�����j�uw�{"����␆���'0��R�������]���1�!IfxR��3��P���c��ED��>c#mI�^7X�������D�V%����������zd��X"��������+,���ƛ<A�U��<@�~�����3��ҟ����zY*L����~��L�p�J��4~@���l�4i�nt:ǪB
\�?mn�eй���Y�p�be��׍"1����I@��20���t.\��_����krpD���3��<3�%����hV�SWFeK�y�䯃�=�S���.�����nT�kk�];?i��-@�'T	~WMEvޓ�uS;�I�V�t9���2��#����b�a�rR����Dʮ;�2�ҌU�u�r��ixzT���S(z<W�@������i�yDߨ�k���5��]ܠ�m~��� ���>3#���BM����B�4�W�d~d�K^��X�R�Nn�F�x�h-��Px���.lU���]V}�SD�b)Q�*�g�%�Ut�:pa(��O�x+��K��8�(R\#�	��~:�nx+�hd�8O�jı��rUEM�W����GNd�&�(G�j�6K_��gV�{��SSn�@�tw��,��J�D�7K	}NO@�!`��t9J!&x�>%$�p�j�)%8Ș�
���n�H\�<�v�4�t�/��7J��?��֒��?q�<V�9��[}����7�{h�k���-��fw�$��3�]IN�A݂6���	���3��z=R��60tWnLY�Ơ&�  �Y�>��xX��O���S�8U��C����\��0.Og��DV�j��	���Bg�{9��rg��g�u�`*�.�Y�Z���e�^���?��M��'�=GY���4���L�����/�)d{���C����B�`����{��M��s����f����^7�$ (�ʺ��2�
9 �����y���@a;���]��WW����u}}��7N�˅ܢޑ�	��T��ܓG�p�X��vș�"�嶆b/���Ӓ��=�^���a��?[�U�q�rO���Y�ڔ}QiV�a��%ݺ85J�:a6e~�t�B�����L[���ayBA<�����s�]��mޅ�����}PP��HHb�#��@[��lȑ��rw\���(�-ک:�n��� ���I��,L�K����X��z٪�)\��'>��*��wp����4;���&^�8�����q�#�۹u�z���X���4�d�͆
e�1DW���/��� H�d�j|3bY�����}_?�<��Ď���mgt�a�����z[�HUB�m_�fn:�R�u� w�*,���@u
�;�d�P6Y����M�.�#�?h���,�J>��`��9dX��)S�^T��U�Jm̬���܌I�Oi��ƣ�eι�O�d�q�KHBl��r�|��	V���3�������M�cxv���_���|bJC�N��Ն�IAWG3�x��Lca�
�S���i�T~��X<����PS��D�l��4rT�*��%�,
O��K��%�v����Qx��w���W�a!I��w�[ e]�t2��EuҸ=�5 _���lC�Į!�'��^%K���]9�*�K��	�E*�f�S�
ZE��x'�NK�Dx�d�Z�F�x�u�Uu�ik� Q$i�sE-�N��W�T���⧙CP�UR+�4)�va=��|�1H��.�ӯ��e6	k+�g9�l�ј,d��q�E��%ꃖei��i1,O3S2����MiWy�F��Ǯ�cؤ�5�{��X),������G�J*f^�H9|m<Pb�w�hr��6P����Zì���r�ҏ�L��4��6?�qҒ"J�u��(k���07ƭ"�e
�-c��ȣefv�F(���E�̉�לu2B��Z%�t��:`�M�w�==�׫�R�z�a[���g�E����������,1�x�C���jс�{�/ܥ�Eh8����Nd�(��	|Iy��ݱ�!�3Dﾑ��H�x�=N��yb!4ҦUK{��Y�0�U�^�g4S�^�y$
~*�E+µc��Gݛ����Q����OS�����ǎd_n����v���W�Uև�m.�<�P���z�O�m��3����wg�c-��3S���X",�1�/{���x9C�x���yŋ���]����#`�"w3}�r�����.-�i�د��q�ų���g��}c>���!ί��/�51һ#,<�;�_d�|so�8^f~��|����]�"rS����7��,F���h=��Mv����2k%�{���:�w�����L�Eu�O��V_���g��h@�3�=8��E�����2��gRr�!2]��������@��s�c&P%����a>.�"��tq�R�}�����i�tx �0^�D�s��c8I�7|�&�!�`)_nA�l�{��\x6�S��яT-[���g�o]�����aȌ���=ѳ������`�����>Έ�p���<	i֧"�"�b��*�>��kX��u8dI�W�Ɓ�|��:�,�U&��g8*;���%x����m壟���5%JP��1M'�NY����$�?3�~٬,RO���� ��9��4��R+`K��;e.�61z"�4����pe=��p�V���'[��K�J��}�-W�﮶� �-<�qGۥԇZ	�tlxE�'�$8�h�\��6H��cG$�;�eMT{6�'G�Vm�{����? ��{N�Y�;�N$�D�����.����b�7����S]~Z_3�BRu�*C��;�U'�Y�M���E��Z��\�Έ���8�C��|�i��2j�g6rq�`،��q�]&���3�o��[���b^s���t�A8񐕸���MQ9��ٗVi�̋��TP	|�i�V�$[�h;)i'^�������4�J�:{�P�!�5(JS��������^m����o�F^(f�k�Nff*��7�"<v��h�����7��}ᆬ��yZ�؜�'l��������v��ғ�/��z�Ac �቉�oA�)�+
4�,�.�ݛ3�h(�/����)Yd{wOL��i�}�h�Yy�ԸU��oz���L�k^�pd�oi��d��w�G����gcX�d����������Q���;�F�[+H<*Vp����upɦ.�Y4)�	X0�`��p�L���t�o��+fz�98�}�-nn�i3�)��x�:�=��c������n�[?ʣXs�eg��9s ��8-�g!�lB�u)������"�>�J��N�UHR���9_��t���w��w���iOo0z�T�Y@���Rm�p�y�2���Or��$��ov�*t=�|&���i]Y~#�U]�;�@s�Ѣ�r�,��u-��y{o|�[3W����/z��'�ԥ�7�b�gI������s����N(�#M�g0o�����s�e6��Ѷ��]R{39#5�;±q�A=�k�t�(�m���x�v�,#6-�jlM�Mx����&�e��{��:��C�S_>*��m�5��*�������/��qS	�yKl�Y�w�Q�>i���j��<*3����AY�f����h^���{z �d;?~��5�ؕ���kU<��j�;����������L�T�'����،���hk�����hRV�ǽ��0"~��Lo�>E�}��i�^ɳ꣜'���w�H�11�0�ȥ\�m����(�.1���}��v^�!��h�@��U�~7�|#a�'z�o7?��l�,l3�EPX�cU8:� dm�s%�j(0[&�����q�g��z*>{R�7N��?�7�۽ɩb�_���[�J��E�Z�L=���j��:\�u��5��*Ug��̸�5��=�/WhO=+v�Ǽ���ԩ����S)G�J�&�G��{�l�K���	�'�P(I������||��4�ncYK��)(��q����R�_'?�6D D\og~T%�c�����̹u�����7�'d�%(��IÖ+)(:)���~�F���^�O��,�����iҶ�C!?z��.��o��k�r'��*s���%8פ*m�t}עOu�U~\֩�H�\�,�A"�>���Kj65u�e}�j�f��k7�n�`�츷�<M?3Ë�{'b��.*�E|�s�˵a����,�Q�gn���:k�5�Ɨ{u`�X���[�F:F�/�f��S<n��+	m���NΕ:V�[ܮ�g�i����h�o��DO�r�.T$b�^�dD�E�4��8�2����h��md����ӓ���Nhx$��a%��~��0��9��т����ۋ��֒��@~?)���Ҍ���9�$IZ���k�L�Bt�ڔq��w��R���$y
�����+]�֛���`.�@���%����{V���ɸݖ��}�F��N��*H5���j�����$=�l��E��a�i �w���r�����+�����,^z���+C��@�֝gH�f�3U:`�s�Ff�2�M��R!g�a�ˑ�m�j����+�4b�,�%^]��3�%�O3��W��̾*�	ݷ�3ВX�೷`.�ۑwj$����:>"�d�c_�2����W�P,���8�����(oI��~�M��*AW�
�K=�b���(����!T&��Yo
�wd�:0��/�v5��A�;�(��b�݂G99/v��"%���f�yds$��|��z�K([��&�gi��y��U��5���IܬG����IDDP�x����;k��`���oS�!8���oW��-O/+�RV�%̪q r�ġz�7�v�!���f��x+[L5t��.Q�ʗ��cZ�.��B�{<#�O�Y��:���ޡ*(����~�7Ix���6�����)��'}��_�L����h��qj�Y�j�p�Ό�4�:�\D�5�i��Ր}��5�;EG֭���|��>��;���K���ޟ	����
�-h1Wf����:��EȰz^����P�i4�qp��E���Z��N�xO�ͬN�ٴ�w�6��:|��3��> ���:���e�� ����26H�C5taߍ�e���Ϫr`�_e���%���\h�Rt62.P��3xfpE���i�ު���N/͹c"�N~j�p��Aj-�f�)��[d���w��aV��U�z����[z��;dWl�EVoZ�a�G�͐@!T�M��@�`íE�-��=;6��1��l\�*���w��on�[m(�t,Ë�ť�ߘg�i�,M̸��gZ�<�m�H�vjY���ޙ4�~�P�cBW���CEH��Z����~�7ß���q���J^o�S,/Y�?��ΜEY��)�E�}�@B�f�J:��z�(�e:Zo���Ҧ�(��	��t�-~��j���߉z�M�1�+e��$����3\�q����(s��-�Q2�r���`����K줉�Ҫ���/������&�O�A��=O�����96����ݚ~��J���~Z0�lf�c����v
|Y_��Ѓ18ז��BD,���4j��ܤ��غ�1�� �(���!ǲ�3:w$Y%�aw�7ͅ�yzf���2����E:9w�6�紛�Q�*�O& �~O�/I Ie���Y��o�rKrM��~Ϧ}�!{������ix����|�sȊ1�ז�6�#C�Vh�^'��"gi���	�H�8Ҹ�^c���@����c���t�(�S�&)�(1��ߪ=l��ۇ)��c2�DQ~����Z��!Ї�rTѬj%�8��2a"��
������ ą\E���v�]�E�q�W_� x����j|3ɵ'��8��	�\����(�8�O&�Vw�|<���e����D-��!�V������AUl&���4s@��?������膇����݃���%T=�B*�6�@u���m���@�X� -��W�a�2�}(����Z��k�gN '�W�H�K������te[�N��KuMc$nۢ~#B�5��!���
��4;�WP6�k�c�.�$ֹ�i50��G$k����wz��:t`���觳X?jh��G�Z���@�ǂQW\�v�"yٽ��o�#�	F�?K����"���;�a�*^8K�4�Z�f�v+p���,�y�|��z\��P	��λV��Yt���.�_M.�D3�1�������O���I'r;;ף߷ ����[P^���X�Bc�o!)��t%맴eh.5��Vӯ&yF���tĔ/?��Q�s���鴃��S)!'em_�������
�@פ{�*�+��'�l�����A�%�LE	�����{[Ҳh$%\	ͽ��γXP��-=Bɦ�,v!�\P�&��!c��8��0�&9���������N�¥�K��H��Φfj�0�6�)�;gD�d* �W��S�i�#�Fؒ0��}�`����[N9eq!�3I�/��Cez�5�LG.�l��B_���|�6r���W�v�����+�O5��3��^�My���[w�A8�Q�hcz)�v�BҝH�I���4;� t��z�����CĦ<&�R\�DKԨ�� om	|`���6�
ć}Tڿ�r���-��x�۸��JMv�S�5��wj���tuKCg��&�� ��6�����m����k[��O4�C6ȧNc��=��,ɋ�b�K9?E�/D[H�Y���2f���EF^�An��sv�D&��G7��.�q���G��hO�,?���i���~�"�%�S�c������IPy���U�I��US/ t�<��,�M?��P�E�����L����Sh�c��q$�[5���H�n�we�/V�	�I��~�2���66S�����)�d���oZ���]�З{?`�t�GQ��&rZ�X���5����V|�<�T �PoE��>��d�.M����Yg����+��9�t��>L0�M�,���Ʉ�q��/�D������mR���'��L:��\m5A�$��ա|�p�\#ę��ԪXGg�xp�A�ț��o���=M{H��V�n.V��|��4>Ga�6�D~'�կv�E{Z�u$��X.5P��ӥ�j��**|V��+�Y�D.��Z9��-_����-�XN$�|�SnY;����˸C��� �'z���br�ag�?������4�v��6�j1�^�iKa�ҪBr�c q5�nHл�!�t^�B�H�œ�+敗�����A�����%�y��� ��/5��V�V��C�(/C��� fD��Lz�L��*7tT���AI7P�a�`Y���0�YN����st��}����O9��},�}b��pA�#�O������6<���G0�N��@�>�S��`,옒rw�M���5�T�la���X_������. ��ޫ܃��!]HI��2z�mX������拥|A��gH'����9FD��\�X5���~��e� &�ۣ�P���P��x�0L%%
p�a���/S�PO�`�O�h��^�b	�9��~׹��jx�U�'k��b��Í�^���)�5b�=�tq� �.N�g��r3���/�u+w����̈́�b�)��K�Y�T��bcM4U�Ü�Dyxf~��nѠ:�z`�ЄŖ��
̲dRkɢ�Ȃ�I��~h�M���F���*�.͝�$���7Loi�xqIh�m�m�ep�S�ot�s����3o�k)����R�y�NJ�Ƃu7�}��������M�K���ȓ��J�(���"�W?*fmp�Y�O~����{ڰ҂������'�9W9�zk��K燉���q�+�G�W�؞N)@����o�d=������(qp������1G�lTX���ĶbLB�F	�͝���/dO덎G���� �K�T�M<pi!����?
"����<v�[�8�~6=!fa+?��^��mB�7�Q�"Y�)�e������]T�LS�|^�-�}����
�22�8����=�`�J���m�s�� J�_�ۥm�#���Cx�e{�B�t�V��6�`�(�5b�������\�	�Y��Dn*�H/���.��o��"&�8z�s�nWR�@�%�ϲz�򍮡r~��Z���5��Æw��=����@��h�gm�ܑ��zlg��Y�:�����|�V��c���݊*\z�~.�`�{7�#�1���t��, z��pX�����<��.5��al�-�	����G4�@�O�l�IZ���πJH���<`ժt��g�m:md�/�Nrz涞+[8ɛ�Y���ٸ���"�SW�i�"�?x'�X�_)������B_<��"��=���uƯ�{ ��(��=�\PE�g pE{�Le�j�;5����W�Iٌ,>��L�W	��K쥉��"�	Q��I7���$��֯/|������:�=��,��ѭ���OU��yP3��#9��@�׍�UrՃ9��T�6= &?���R͹?�[Z���G5S$ƜIU2��xSZ9�&�(��HHe��o ,��WO��X*�!��������zJYTi����M���3�K,8j���"ȞL~�ATgU��J��h1�t&�:p��cp��u"Ӊғ��N��ѽ�6Ҳ��efq'Is������-LM~���ALXF�����N�i'A>�y^���#7�Ч�D�
�C�T�@��fl�dhP^>tw�f��\�S��#���9YIa�~>����C�.�� :�wt�cQ��5��ر�Pa�$��{n~RX�)�.F#j����n���[-屁Aqz:����X�*V���坅�#���^�j�s1���g)��t~��N�Ę`�k�y�I9��Wf���x�]Hh]�Eг����,Yg�^���C�����칱�б�z�3�A��[~��k5�f;�O�7�W�Z��/�l����>aD�������pK��b���;���@n�:~ma�͛�11`"��˔�צo� A}��p��J^��Q�F�YL��]���6��4�"%�&��"ٖ�����)NFQ�Q����3qߓƖjK(�-� �V)F�9�t�d��]dt"a0���ܒ[�#������ZkQ[���6Cb	��L��3�YY5����KH�;��z���i����3���.}u'VV/�d�+fe:�T����֍�kݺ��y�&�������v�-=�p��Խ,����QCG���4"�n� �C�A���V�8�6K:�_��+��=�k˥�R̿�x'�f������h	�@rô�,Z�r�0;=Og|��O��J^���=���.X��PD*C@��IB\b ��?�s�F�s�?��I��f�OO��IO������o˱��&'�E�6+h.U�4��wU�t���k��?���":ȧ<�X��T{�	��3�~��r�/��7\��I�q6�g��=b����d4z�g�{}���ꛛ�C�o�v�ߔ����j|㶘�3z�B܊��\)�*�1��\:o!/p�z���3�3<������:�J�.�9X�yO2x��ox �7y�N�G�s7ܕ�����F�k����4 ��pa%�Ĉaߟ����8dO��'���Zm��g�����^
�C�"�����ݴ6W��o�`��k�kgt�#F���dc;�<��'�qꁀ!.C�ݻ��V����$�U���-GD��F��!�vԢ�|e�A$`���VWɮ�C\M��9t�/	݅�5<h�z|�0�1%"��Ӫ��R�HǨ�+�"_�ݖ�K��BW}�[N�/��U$�a�f���B� �u�X�IK��Ã��u�Q��9�RH�Ô���6BUݕ�W������b{n��/�;0��d+f=�&��:����#O�$U�����`�;���::�p�޳�������d���24�9#�r��Ϯ�:����r�\��_!�)Ą�G0\݋�kW�4??�K V)�B��p+*lj��գ"̭ylml�30!h�]1ۘ�]��>�����X�zX/р��S?BT����;�Ή1U��`TBu>3B���.�:����?�I'M'X�[���ڐμ2t��%�kϛ��a��4r�_ ��د��n�ˉ��q۲�3޻�b��Id��#��P�!��rjz��c��<>1����~����V{�kqdV��
�'<O��yw����W�	�\ͬϢ�Q���|��m�(��t	�L�4Y�pʳ������e�'�c!ٻl���g������*�>���=/��eA� UZ�b�Z�ۼ�ˁ����X_���6V(��i r��O���Iב	���t�J\Xjk�P�2�D��qN���\tm��}L~�`P���r�n�vZyi�;��g g!?Cs�o!���1�,�M���+TC_W"p ��	�Y�kBJugs2��6y�N`�HF{?�OBZS,("$���<�q��]%4�)8���<�+y�qr��/Ur���BS�����]�mdECci�8P�tp@5b�0��T�6����4������?G8�߆9&?���b$��~��wG�^�)���U&��1�\Q�t�R�+�P��ؽpm��sXie�j{�_�n���P�et)�E�*�tO�H������1zH�,T
(&gj�����UOY|6�@!�������T#\x�A��+���"n%���l��<bM&q�&D�Él�N~�TB�#'͐6���-����|�A�̡)�t�� �k(���kW�cNDOT��˝=�l)��@�`P#����b��Ͻ|�2ͷ�2t��X�p�������̽�u���L��T��A�%_8����w=�k�J:��y�ZV�g�]/l��9�V�Ε�Q�̢����F]�_�7�z����-$�4g��\���a�㧛��!$�>F��W�6M��<��1P}x�c��9�K��θ*��dx+�*s?�t���j��$��	T0��j�ɯ�F�m�/��[hQ18���d�������L���N�5��'��F�F;൧��`S���ʁ�^m#�8�k�0��H���Y���%�M���B��QjR��4�hK6;�#=��<�"Q#m�s���]�1^n��g�)ĥ�#j=�.:��R���שp��=��`�2���>�ܭxٸ����_��G�5��@��0���HnO_����ԩh �6���X?ڤ`�q �j�׬+Vve�(���?i�}$0��d�'S�t^�g7!Y�w�jHE� N.q�L�1��� �V�w�dF��\-�H͗ׅ�g�BA�_�þ�(��#����zC��)�hɁ�U�M������C���gd|
�w/v0ܜIָ�a�zg�:�����䲘B�%�#^m]C?�4k�1�?����.�3S��a�!ɬ�6��H�&�y�,��6J��#^; ��E���&�b�e^ی�Uw�ûD� W���]��4y��Q��L{ĵ��ᜓ�<3�U�H\���24�TQ���w��N�BF`|^��!�1��d0��'��C���0^�'̔W� ���
}�������Ξv��me��!,w�C������ax�E�7q��W暊���7bC��jP��OG��m���7���uO[�
�V�Ж�F�ߺ�&�.vHt6ӧW���]R�S�¬����S�9���.c�%��<T��{/�}W��F���v�dB�l�Oˮ�un�k�e�a�Л(��Ҍ%�]�^N�z��<JĨ��")� ��.�u��7f�nP��pmK�n��{f��0��E?L�N�! k�)���T�S���Ŗ)sä��7�����8ʍ������7��Ԯ�f��i��C����F��b诧%M��cb 䥳T��
��ׂ���EHTӉ-6_������=�v#�����ߩF�)z{��TКW3�tE��Th���g�+Bْ�и�m /�A��~�N�S(�k�7��f�iWA��g�=pQ5�ٯ���� ��.,�A��${}�%�J��=��k��ȅ֌�1U�Yl2f���ĿY��
P�k�9�"�9o��
��L���tw��� ��M%Ʋ8�G.2�5K�%�5%oЌ�	��oh'Й�a�<�[;�|��d��N?�79�藝ݦ��v�9��Hъ�H|=[�k�@ S�xaE�K'�c4V��-h��"��f$Q�J��A�����L�C�y�\����}qC,m�԰\@��/�� ��L�Xk�|�0���3m�Z�������U�
ǩ���R֚���>�5;aؤ7v��=sN��hx���e1Bvz��O���F��ɫ�� ��Eӆ$T�N�zCbK{U�2+��ѣ�1�lQCd�θ�<󉕊� ŀ��*��+v�a�o��&
P��8��^L?����}
�	�Ȉ��^_��4YNA�(��}����K����7m�3��?zw�5�rw��f�����JG��^����:��cY>i�P��>�5v&�,���I9�>T�{@�}U�B��K�L>U��FkD�x�j�r����mݢ���$�P�ޅ�E�e��#�?���#��1u���[2V#��XB�N�i�_/%� G����D ��괚�{��&��Ar�X�3�%��ќ�0m�jp�lD@C������~�^��Y��Qi���	z�nh�O2��<����8�~��g�N�5LT1S��H�Y ��Y�������~o�,������4y��ք" �熭�l֫3O�U������M�{r��Q$x2�B��5Ϗw�ș��!���B�V[<����L�,��j-$*�~�|�O`�к�R����]�� ����4h|�d�kS$����'L,��9���휙f�Ia�g�D��`�A��#�$]TE����6�M>�����{Xhft�~������7���+�b8��x`>,ݕWӮ��@���F��(Qz�V�ՄN�����Z����[KgB��1Avo�ZO����^�įE����,�?�y�a��]�X<��I]T��� ����7������2\��JE�<%QH_�4�(ܧ!��X��Vɾ~]��6,�ܴݝ��C�P�%Ժ�W�۷���BJ4�C��?6վQ�����m�u�~m���՛H}�q��`���3``��Àp@T܋��'��#?'���jD����<�����}]��'&N�VHfj��x��->C�.��J�I'�e���Ǟ�^pQ��%�a���r�sh
M��Սp���1X�J=�w�l��ik
���ޅ�i�F9��M����yc�wP�;���oKh#�/�W%�r����q���W⸠�Ƴ�B�?a��l���8I���;�Ai��k�8��֬��1�mXA�8����X��@%���[y�t�j��R
�����.��oS��4�K��5�ѷ���O�1�i+Fh��� �u��ۄ�N;�їQ�V^�
R#����a3�n�׏�"�s�wCBۜY����y���`Ij��=�_�����Z'h�����b$`�d���g86L�2�����|�]Co�TB�i�^.�f��bv�q4<�J�`f��I#���]�zYpIAF|��� Pg�����x��7���s�3��="F�`p���NhEWc�u��M������l��[�>��Y��OS� ����h�0y?Y����R����5!n��飽P�H�4�=�f3�s=������bP�^%i�7J��l�c�NĐ�6�k4Tp�~��²gm������m����3�4�Rļ�5&e��1T�J �̢@���+�Po2>
�e�K���O�4�?��|�m8� ���*B5�j�8�Yg����q����h����k��߇�Cm�{������0�9�Wj
↭�.O*T: �}�2�|�(�k	�v�?
���pE�>���@�*{��[GTY\�Ϭ6*���a���s5~J�/��k�h?���igV�m�}1b�B����G�f�uE�Ya��I�Ʊ8�$6Z���e��њ�Y�Oȟ�^�m��.&�Rn@��-����&�?п���|Dn�1e�N��Sޜ�h	�W��d3�e{���L��8��ǤQ����	������?!_��\�W�(�p������c���W
��T@Qj)8��7��}� 2���)���d�^��F�ŲB0���|B�i/k!g����n%�~]d���S�T]�n��2�>O�eD� ���)in���Ѫ�$���c����h�TМ�ۣ2Ƭɶ�@fq�Y�vIt�-�Γq@�2_}ϵ��e,�}�j8 �Ī�m�LL������7�ԎT���?�5^;�Rwkt�d�V�Lr}�������?�%ۤh�FF���:i�!<��2����n=��ti�@J�^��-��.c>���X���`��h�Ԉn_e����\���Yx�����̵�a�<+@���6�����b9�����	v�<Je�u)�Y ��@�&Ӟ6�D|���������2���NONۧ�p7d7�)mS"���oc�j}o��M�νmj�������w���m_�f!�LOӦa�P�Ҁ!�HGԆ�&�����a � a��{�]{�~�(Ւ��Y��X<@ �:���D����0k�8C�w�J
-n�D4��y`�8+a�[//�M�-e�q��G]҃��s�$�f�Z���,5݊ϙF(�J���ˠv���)B�\��R��І_�a�`mC^Ӝf��m��.�P����H�ei�'��!��)٥��2�CѴXx�%Ω0R3}�@:6�ΚOn B�(�8ncXw1	#�S�<���A��F����i!�ȕ����{�V���k������=(��>����tJ��гU�-�5�
g�0�i���Ϸu�M���&�*��7�����S�%�"�� ��/�{�����A��Q4�׏�&½���xcRK%s$� _g0q���n ��(`:n�&��C0V��	�x����r�R�f��w'� �)�o �v^l�Q�"c~c�hv
�T��P��: }E��.��9�#x�RZ�*���7g�\�X'�2���JK�މ;te���Q����c��2�2vz��u��/Ǹ;gr����?���	Hpn�@�?����'�Y�z;�p˛�[ㄽ0��Y�h*/�L���l�<}���:��VI���5~�?�c�!����2�H���GRH�;'��1��%v�MzwZlZ�gc;��"���`_:�?��"ӣ
��ǰ��D�UQx�	]à��j[�E�_���<��� ��  �����~�y��(4�ex�=�_�>m0h�ߕ�+��܈�O�T$�k��RyKYB�s,�r�G �M9���޻��z�HA�w-Y$�]�E0�A@G�����d���n�V��H��R�_0t�9g��d5D�D0^�&d�9x�&w���(�`��֑rN_E�Rۿ,bBT0�o�b̨��'�_���g�w�Ùӗ�!�j�5��ݗ��/���T�NI��0Q��ǎJ��I�4�bZ����C4ĵ�L��`���'�fBH�	*�vk~n�ӿ:�:`��y�g����=��l�sa��b�&�{u��6�%��jn}*N�2�t�ބ��6;	YQ��Ͷ}e�59���6`1a\`y�	�3�.�dڴMj�NFX�d�LAT7YF̍G�VK*���MŃ���D��_�.�c�dQB"{�����+�Q�P&�\�?2K��`Q�[�/�<*cJ����oM�*?�T׎pT����P"15ss��k�y��~����w��� ��aQ���V���nX��*s$Ds�u��ɠ|�8��Yr�+��0�W�3�x�;�Q|�.�1B��2ؖj����[��F������fc�o��U���TsS�<ƒ{�������/�	ˡ#F�6��&���Wa�r��sٶ#��E��-�+U�N���g�Oa�zt��EE Q��4˳��G�t���[�`��$L1�b?��w�璓~ȏ�Y��=9�)P�&�җ�D��"��\� Y@��aO��%���6៯���|t8G���q�Z��XL���s����1�c �k���?.Ƴ�T��	G�:د4�y���in/~���C;�;�7��?������K�-����:m�B/'��K�s��7�S)w�1�"`����!+�Z[
AL.���@(�Y��-ӵ-���v�'H�͎>�m��`�k�s�̂P���F���J~��@e�ČxUH쮪�'��}4�^�D����Id�OClq���^�ɹ���%X��a{����jR;:��V�n��q��F]�3M�)��v�b)Q+���,�-Q�e�
�sf'|L�E؇*b`s����V�����QU�������l���AZmUuU���o����)��m8��	����v6O&�L���"��l1ʛȊ���rswy�m�E�l\���W��w��4�˾�_�ow��vz�_�,<�%�������w��Z���Q~�ǵ^�ڭ;��0�F�U7���X�B\�5ɜٝ1���C������`���`�U�<�L!>��i+*[i��Q�̜+����J�ۿ4��YK7׻�^�a_@�S|�'��p��N���08�H#yK�,�6�+����}3j�OZRd��ýBf1�9�IJ$��×��>X�z뚒=+�	�7$:�!���u�'�c��%��(����qƷ!��NA���Kn%� �3���,_E��"�W��w˔��=�����p�Pd9�X�0i��\ӛ�mD�WD9�΃+�?4s\~�?���n�' ���Z��~aa�`�=�Z��yw���+|�/iUC�,��sxL�	+��)D1J��,C�L�{��2����o��5�p��^�I��g܌�����ie�����O����n����E��."��sjhM?gR�3�L��Ï�q>�ċƔ(5j�9N��eK\S��m9�+�I�[j�I4�ֈ�I��bp)�:��8�����l�j��Z�<g����F��v%�(PS5дk�#��_2���/�������aQs9�HЗ�:���S����R��
M������
�f�(�8��*ލB��gU�)�]��tח~����0g6�pO��R�U�+��4Z�M|S��(�o =f-�S����ڵix�����^a�Ú�� +- �ڶ-��7�n��	,(�5Sm��u��ګ�<Dp��T(e2�.��y��N��8�C�Z8�d�E �p�M�����+�:y�����.�M��)w��#�<K}c|��X!���99!��(�ޮK,��w�?\�6֕9�xM���V�k	!;j�E]�ud��"�����ᵀoY|Ӈ�Ʊ��aa��c�Bv�>%>
�c��p5���fƥ`�d8L�G�se-w魎���݈�@�!�?Bd�9W�V���x���wKݸ"?^Y����4������!W��8���X����X��g�ٚ�62�����C2W�1��=���=��
 �_��E���p��j�bǢ�$;�{h\�W?�3l>ɵ8*+�|5o#�0~��[�����ƺ4Dd���1'�,�%�?3N;v���TYYQ��z��Q��B�V=�?�<&6@!����&؍v�oA%	b��" XF�6&��\K����w��>r�vWJ�[�xj��1Jh��4����G/���e[Z������&��:��;Ca[��]�-ݬ'�JÅ�/��.
�d��c43����:Q꓾�h|�B���ŧ;B��Y�Ъ{�'��c�� �)1�͹+���͍����O�����}�O�� N�0hJ��
����b>�򃳡:���#�>������q��O�M�O�����|�ϛ�I�醴��//!G�gd�V��Xm��k�N�j��`Dd��H�7-�g+�L8i�b,0���z����d*���&W���Q���.r̬��o7We������D1[}X >H�:��gG�/(����}�15��1�#�����+�>G��W�#� %'�)�j]�!����N������W��ٿ��ն�{=g^��xfL;;!��jY4o�C')�Y)��$�5����L�z�E&�?����G"Z� U4{� ���M��b��|�^��vT���=UÝU�nrv�!9I��"M�.�sp���K���b�,���5��'��h�7P��#N鱫����%E.^��y��%���P�ֱ�RS{�������zby��"e�]p�7sW.-+�.k3���\Dm~v �b�x�z>�~��ee������<��0Gح�E6��,�#n��g��Ar�������rQ���Z�����Ӥ�T|W��C�����/~U�ֳ��ΠP\��dA���>��ch��^��W%��P*�]-ń���#�"�]h�V�|���8�����h���t����Vᖸ�́�-�6܉�ܝ�1��J�X{�3� ǟA��F������%����`�����R��kZ �ى��Wp^S���I�h�#6W��Ė����ҿ#��Y)v�_�)Ҝ2Az�]�k����Z����}�)��J$4�^��S�����'��ܗ��Dжpȴi6����iq<k�����v�r��[��B�/h��+�]�9vBQ�!6����OP�d�M��1�.H-�Z���INݯ���*Σ�gT�nZ�q���H֌��m����ٔ��/�D-jFF�0��B��51�s���:՞ �9BN���`��cA~���'#����S2K���qjp�2��6�Z���3W���� z��4� ��ui���DdP��q�l��ݪ�=��g��U�KE�������e�0�qF��릻�O�W�Z�s$ː�|~&ty�Yji��[��bf�*�n/_�
r��Pd ���V��y
4��9���[<�����Yl{F-��aN��
DjTk�~S�vj�M�o�' ��e�i�gભj��eP!��]#�Ю���?��3�u�����8�vI��/y�:�^rQ��=� �G�V���fϠ}�6P����7��ct�UP�3��-.V��,{'�ѳD�Pa�w[{ʌR���������$�9U��S������Z<M��-CpO��6+�(=ѫ��l7�T�'ѕ�v��O&�D"QV�.۴��T*P�]q��{w�8F��w�T��;Yԇ��v�k���䥠�+Jg�5LZx���踍�&�^���X�淐;p��YfyUM�9��n캙U�t���O�͡���Y�KGe��k��x�ۤ�� T{���Cғ�������NpȰw��-���ъ�i��cP���U�a��{��,���-���̬ԁm}bP�\(9*�N��{^���D=�}c��ϭ�fi}t|��)�kڛ��[~����f.��I����<�8���A;q��tߜ��)W(\f�x�V� �J?�����4� ��ӖZ����N���'_f�o���{����~�v臨�K<B`���;C���'L��o����]�b$�ʆi'귷��W^�Eۍ�4�b�㑛 J؜����u!�{��ʟf�/$�H��٨\�$��/��7�tnp�S��4>"��yʐ)6�1��h@��c<0���W����ҙ"<\ywf�(�0�ȜDo½�+�>9���6��'��p*r��b�8���3%*�4zy�>��t��8<��4hU�
0���P�Y��?X�z�=p�A�[�i�<��ܮWU���:5� GФZ9v*��'j�/��@!�]�1�Bc+�:�l�9�\v��(e~ߔj/����֚4ݷ��<�g��Y����]�~��n�~f�
�Uq�	����:lG�j#����A-͡��:�D-+o���<b�k4�_a`V ��֔�����8q��<|��
rUX��.<�_+z 8$a���꤇םXW�z�
\q�v\�P��q:}
�[2+�!�r �C���`��&�F!q��D��g^N��}����-}�K����͝�|U�K:�lb*	��4جa��ХV�r몠�����~����zL��-E�8Y����(�R�0G$ߢ;�����zүd�G�����U(�t�����q�M"Usk��=�JP�.
r�~{�Ynd��?�2��X6��N@��߻KǤ	{_�ê���+�l�r��b�`���k������1ą�/4u�pZ'ק�jѸ\P�t��[x
o%R\��;[����N~<|��u?�^�ý?-f|�N�aLL�������ښ�keڇ� K�`�W�rc������K�9J�G(�͹ᅴ�W����Ts)R�]��J�fkI5�@�/�V+l�W=;�mdAa���=���K��:���2����yZOfV��ç�]Y��t��o[#ʴ̀����1$3_�75��P&��z��5�Ճrw E���  9���(]��|���⡜��r]��D�B��
~	���6��aQN��<�R�AL "��'~�J��g(��2c��b�p���2N�r���C�0ʘ�Jޞrqs���{���q,�؍x�����ao�vYʪ�o/�+/�P�E�ǎ�}+������Ar�#Y>��؛��ܐ!�d5�*�i·!帼X��p��'�}1D.h�˻�fm��N� 4�0����%p�^B
]/���ZX����LBLS\b���hF8�'%�"j4 �$�qte#g|�A������~��2g{�lH{�Л�A���M>�������_�yv�IbP�o��E��%�˖>�'����ĂF"ɫW����4{GR���VoFcI)���.��6���,u��_����A3�&�'���0�y�  5Am�i�(��sN�P�n�̺��Z��O����)gj����є��d8��"�@��<����ڱv�Kƫ'�+��MAT$��t%�쨝1M�;�� �_�-���3����n܃^�m��Ħ_c�+��w��s	���;�6�r�!���fT�K��:p2������LaPԬ���.n�ì��7� +�Z��&��+}&]�h�b�+���T@����uY6\��(z�E�D���8އ�UIء ;J�b]���I��N�w-�u�C�S�CM��3~Q�z̜5���<[�E�0y�i���,=�c#|�
n��W���ˉ�m�9�aO��vr�7�_tZ	Q&��_H��>K�u�&&]�)�*cA"H}[�QZ��,Z][�z�KI����:���Ln*����Vj�HS�<L�/=��-��D5[�"/���Sx�b��K)5�%�R�ř�hްJ��;ZT���7�kpn�V�$lEs�Ҟ�d7�?<b`�g��y�F�$����Weu����յ�m
��2	A���M%6�a憬�23ү5�՛�P��U��l��w��7
u�w�OK�H��̚U)a��DPǴKGK�wjI���"*o")��rK�X��������>4�P���C�AJ�+�FғƕJ?&/q��:�52�-oK���b��p��m�@K\D����^�ĹS˔Z��	��p�9֣u�����({)ڍ:�e� �^5���1�nl�"���"���6��ȫ���.@$�o�o���JͶ�S�<X����LǪ|����.7Z�
W�ݚ9�s���P��� ��⚢�'��*��2�9�E�<?��C�K��9Vմ��{��.p#.�,F,q0�� 拾u�2�v��6�Q�7o6���Xa_L���Q�7)(ޮ�J��P��f���iX�[F\���O �jэ]͏:��Vܧ^�۴���|Dz���p�~UR�e��li���h�.��x)��Z�A����ղ\��Y���ߋ3��������V����a_�o|�L� ��l�Q�ӌq!g�]�7x���7i=]�iq��>���+ގ��|��T$�|mY�ߝ`5�͇!�j�.�i_��L��Q���%�~w��_���D�l��q2��Z!L;Sr�W����B@v�4G�d2hxM9q��ξ�&�R��nݫ+��][�&d;�1�3��L۱�qD�\�5��_��{Z��U_=b���H-D̻��MW�6T���t���ǔ�O�4g�"k_ �v�q��ƕ�A�׹�肂���S��ݴ A���Ǳ��"��A��ׁw�:��#g��6s��=�<�4$&U�&��� CL���)�)�pe#�~C�����o;i�)���76����gUJ�7����	y7��w*�~g)7d����������]��F�����9q������5s��O�E�\-b�!L� -�5%���Ţ��9�ԇ�*~��p����x�4'<*fx%�1�5L;T��O-*B��"���I4��R��U���bϋ�bp���
����0��������|�Y����o�E�.�{�BAəB�/*���MN=&��b=/c�sOksfx�o�ֹ���� s���V~i��CVq����5=Wu�R}�j�	�b��4{Z<r�ek��ŝ ��gdr��E��|�8�?�ފ��K'�A��@�m�����P*��L.���'�����a��*ą �K�
�����f�ܞM���aKe:�ؐ3�@&�V}� `�Ŏ��������D<̂���{�`ʰL.�0��X~��^�I����U�^A�-�_�� ��HǬ�s�;9��(��$h��&j����=�-�>�u���n�G�j�L] (�����8����ɬ�{pU�G����RJ�yM��av�U�R�1�*�>Mم �y�?:*J
��=�`�Q�ɮJ��b3羝������o��g��րz��i���-����h[�U����"��o|�]L��Lz�Б6̋��_��U�w����@�@���
\I@(��,�����ɀ�:o������u�' 7^dk�{�:i���-ɻ4���\��k��>���],?����H0C�:5pfQ�P���ը�׍7��m7p�^2�9�g�F]����������Pv�����TT�H��j�n���輝�EqM��K&L��	��+���Ѓ�.<�����{���>G� ����<C��Z)F��q�4�����7��?m���7�ӓ�?LW������*�qK�����E�����<CᒦK��&�(
تgL�_�M���"�7f���AY�a@���Ud%���},��r
�_��u��υk���O��w�	W8���.q,��~�x$�PK�'���+�='�=�j�f�f�����\�[/ʢt��G �#_��
V��N�77�w��A`��:FI��Â�ͯ/�b���+�་�����SȄ`�J�-�������4ړSB�0��� EQ"�X��&��b�p[�0��������E��GGP�����
�.a*a-��-s\ǯ�|����פK��\�в$�*P���F��f�6��+�4=�N��PuK�φ�pv��I<��||��*�rq�	�gw��&n5�[�`uv��1g�X�{' ���(�v��/��ݍ<�{	m22��gv������%�ț�iDF��e��}ô!�1ڃ�:���5�OG�-�m�f�
?Xn�ֹ��
36B�z�fY��Bu/���R?�Ţ=�x�k�!e�ԃ(�zP �=���;�����6��(��V�n����8��	�u���)��k�t�(��*[\1�y�[24��jܮeeC�ݕt�Κ�쵔�����`''h/5�Ԙ250�n�ﲤXJ�A���wx�`T;�� w��+k��w���ł'��#�T�iT1.l���kYGz�>2u�s	�À���n��9��������*��W�r�{�g{��3P��s���|ƃċ���/ف�g��<`n^���{'d''�I?`��d���e��<;��0-���6%NJ��n�����yh�Ć�'��������Sf0G�#�Č1�����]~�w�)7�t�(u��'4A�OuE�	���d���Q5"���9vh� �YmT��������A�nR�z`�\�!I�s��0FC&���h_���;9n���wHP�YHq�0��ִZ�!��wz��fҸ�4JX)�#��Y/o(��T�+=�͓�䐀�
�N2!��uT�O*�S���1�6jfiGq�gS��[y�
�%"�e�C#��w�9���X��t��Z���;�j��0|ȑ:������b1��+2�Lh7�%��l�琬�=�7�x�.^��d����P�c	m�����v�Z�C�O`�l W-0m���v�͔�5t��U(߸�G�r��5���Get$�:�ͼ�k]�/zC��=(�8C>��v+�yO#�7撪�6&�`Ӓt&m3;���6����|�_�-s�O��n+|3���@%�-�������`��2���q�Kݧ0+�P�r*	 ���'�T�°Q�sӮ�rEl���5�$x=�;bܿ?��"��_*��'���Z��N�4���$�zf�x��#��Č���X�z/��y�E���#��6. ��Y��ð����
{.�Z�U5!�WI^U�&PA��rX�v[k�����v�Ӌ�w�E�IP~�,��O,�nWdV�� V��ZJ)=�F:��̥�|L���LDB������-�9��co���|&���m�*�m�kG���8 ��g�-P�djN���j�
tB�Cl����!Iɴ.b����@���/H|�¥)*C�*���9_�Tq�w������g�W�`��Tz��`�(�|��ƍ�T�e^���x�h}�������>�hJ����2k��t�nFE7����n��gY�\�ϰ-
b���_�>z�I^��q���35bhO?ÿ	Aj}�(3k%c���h�^�kdl�_�?�ti��Pf�D��q����Co2�ɰc�`���P(?
=��8�V���׺d��*�kcb�����J
��h��ˎ��pg�C&�Y3X�\p�ɹ#?�QUg�����{q�U̻Dr��zZv��̅h�c�f��8Q���f��xk��U��ꖞ\P�pk;��c�8\|�&![�볞�p�	U9�k�)��MJ��3��Y�Ӵ��5��MG�䁆8��E��dh��� �,��!�E�t�/j?8�� Rm�����j��g2ظ�ե�,��hRb����G >�����o��[�����Oxxm��h�i���!���Wy\�������(t��}/���oo����<̞ �X���o�������,B�'Y-�J���m�tv�n�[�����D9���8��]-뷦&uqP	8I�c���z��٧IT�/����vewI���#3�̄�)��a�m�,��}�a�̒:q����l�_�؋I�N�w��)d0e���:Y�wj�t�~AK)J1�
F��9�JGҏF_B�Ua�K�^�cS�AfvF��7� k~��bFyUh��IKۧ�#�Xv�k�4@��i.�m�.�/�e]2DJ�`!�u���ɫ�U�� ��^?�_��|�6M]�J�]!F	䓪�U�Aυ��$CQӳ_�)R0�궘��7���������k7�!�Tt_+p�Wu��]
dF\�;��;i:GNzi-��d{�� ���1��@�������O���㣖���`�]U �WN'�����xb��R���C�c��lSDݽ�I�<���#���p�	�,G��#��f���C���{E�	Y^Mb��Ks�Őd������~�1(n �'D��󦍼�PX.DI�h��$'z9�ۧ26k�	`SJb:mnNS��@�FC������*{dؿ���=�:F��r���`���Y�p��hmy�C�Ժ}���HR�޿�"�����W���ծ��"�Xw�v��t�r�A�!~��h�&��K� ꗛ���Oe��?��Q��`���������s��+%!��W�D����h@-�*�zF��)%�	�$��ZD�4��݉M$C	�5Q��D��`�<�[e�v��	��]�;=�O����c����n1�6� ��6@)�[S-n�_�65`��'�A[�23��t�*��r��(��G���\ߩ��1Ϙ�9������m#��B�06���K�L��w�VL�ܛ%���l�C��n��?
ШU�U�;�<ٺVS��lp�^����y������h����Yp� Gx-3!��׬oK/�;i������Á����V�Z�ϸpeι�� o�B50aZ-�n�a�Y�f4��z�Şu��N�9�8#I�1�V��ű�=�%���1�ܑ�}��1��5�)sy�S�u8�eU!g�:KkJH�@������B�A�E@6��IuX��6T�ǂ����\�~=������W��2<�!"�<�)��6��8�[���6��{6My���3��6З>��WQ��A�tt:��WA�x㪘��"i�&i���y�+d��ӛ.>��U	��/T��"�ґ>&?XF�0�Uv�LH1S��%h�'�sªpX@�K��~�	�M�E�]���`&�:S\�r由��]q\�������xc8�XK����ҥ��hA���r=���^P�~yq���,���~w�~���Iz��-
*�وn����!
(�J�ޞ�.@�IoLܲ�B�x�-oɢ\/|xB�ك���/���Q~ Oen� ��!�S�3D�b2V�5�����x��8�#��ʰћ�ϲ�&!�������^��B�7��*C��C�j�]BMU��?��B�:��ʊ&g���N��T����Lv�^�tϥFy�ŵ�|�6���+C��P��.P��;X�u>>۷��%R�05�d�O�o�\��ˈ���3�J���?M��v%��L��]N}�ǣ�Dm*���bD>�n��ln���F�`k0�����ݠ�tE��gw�Л�P�<� ���[�%����E\A�˥-�f��/������W䢑�P�'�4�3kb��"�N���T1�hj�;l�|z����Ȳ%�U�bq�����`-�R�F�񞤨���/c��bl�1;�E��]�ɼ[��Iors��>�S.(��zkm��誦��Xv(�|5��� �[O3��^�uR@qH�4�J�r1V�z�ؒ��$���jh��9���%�`�e)!��z~�X��s�#�x�}�� ���]�ƥh���oI�#կI��r�N��_�Y�1��	���2`�]��޸�F���hE�Y�$Q�.����:~��7�H\a����.η����\^�B�5q�2;P� �'NPX��Q}z��2�akx�$�/m�b��J}�"y��\<�J�+����~)�\띭VY1R�����j��E��`��FQ<��OvN"�C�0�ʪsNq�ࣀl�j�d��$v�9y�����H��!:Ȳt��tE�x��\ܰ�}�ܧ�?{	߮�
�sURĈ'�����v⸬,/��x�6E���nb�Bw}�9�o
�`5y�i��uq�*��?/�a�;�K�W,:g�'0�K�� ��ih���U�[b��h.)a��k�칍�j�;��Ŏ=;{������H�
�h����BUȆ��7U��{v��s,e�� f-�
�'O~6.�R!��:�xE��Q�/s��K:Y�8��e<�x��Nq�|x�����_�Z;��=Ng+ +�7~7�`Mj:␸���� ��~b}��:�`�^��"��h�4̇U�ly��2䗨��>t��w��/���yY������
=�׸jt�o^dq �S՚��R
�v�G��b\�#Jk�qܡ @5�X#��m�����������u��S�n��@�EE��8�5����b�C�!s�Az�ѼW��vq�gH�������
��7�±܀��-z��,���'�[�h&�*R�
�c�6 ��8#��2.�E�y���pTr�>�$��\+Uz�t� {�*CR�V�*_4��o��尩>FGR�} =J;\��⎈J��FO�v�#� r2\;7�q�9�@�$��˕�����k	
��J�� 'nk5+��q�
goF��Ho��7��o�.2���˟a&b���^�f�%��Y�g89Xw� ~�@�Hb���XC���"��?���2�(���#��H�e}9�Ʀ�X�G� ��
D�-*�I��	����W�-	P
�����$]��X� Ѻ~�g�|G�#���zTTm���@�|d��[�ҭ�ch�/�m%��y?.x�K4�v;1�l�������M�����1s��+�}4���2�s��Z��v$��4Ԟ!H���gxk�
��i*Ny�`="YԴ:<�:"�:���x�>;(�"�;�J?�1�I��G��b鎦Шb��� 7���ь}y!Pc��)3�*!qSC�� �d\X/l��8�����P$̈S�UUZ;�߲�wЀ �f���F�=�b�J��P��1͋t)�S��D�?���䀭��Ț�{N�I�9Rm1M#F�CwW:@0χ�8�>���%$9l�
��+3� �|��F
ѕ�i<�<,~g���L9��c��:��b�tzS�b�Rc�����v�{/S�~�~ƍ��F�_N(�U)��St?���9B"q�h ��e����7�+�-������LEХ����c�J�n Y)s&;J;l�M��ٺ�6s�O�A�q�ffi���^~�h鯬�$�x-(�b��/N�9ւ���{u���_��e�=�f/d���P�N�חE!��8k�/P��<���ܭ��r H>�x�k^�d8�F�;�����k����{�l}p��H�S�ʉ	���+ *�-F�c��þ�M�3O�Q����IR��X���p�Ic���tZ0��5KN���; �N�;���U��''�ۜ��}����y&�C�
vt�9h=��䝠.e�M��'�2�m�;����<e��A��"Y��g��ϧ�B��3��
�<)?��-�֫`�����4DQ�咨?����Bm�默[?l�lC���u9J��-TWK#�W��0�#K�d�ɫ���J���6Z`�q��IS�f<�P��!ٚS��`3l`.��L�&����a�~���5j9Ú�D��b-ۉ�H�FG����2��.ϖB��0d�T0��{�*b�|W��^�!�p���1^3�I~+���gۄ��7�h�D ����9����
�>����eөXc^���\�����2 �ZCj��,h�2������up�DO�L����Cr��'�Y��\��ޅ��g����a�;ǎ���1� ���BH
؆Wt�
J��z���8�P��2����,�j(�#�D��lIc8�M�?Xw��2��4gW���Nj�9�%nb6��(����^�	�P@���>��=!�i�v»T��!h�&ND�vW邗U;�q��ܑU��{�"���}k���7�6PB�n���m���8)z~��	��b��f�&��������L:3Ʀ�HY+m��/�j�w���J���#XF�:g�����3)�Ff�S@������rO
�:�8�������� ��k�a�D���.���}�,����7��:T#�
�\��Ip�J)K���G
X�d�L��dF��wS2F�����n3�8tC��rO�w_�������p��"+������nG��@�Z?��i�⍊�<g��=�:U4����E&K}&n�A�XQ����a�U��t�'��>��G<n�O����֨��8N����W)K�)���c�N����Ru*�� 0r���>l��j���\�y����=�������#������F	i�h�~�^])K?H$�����I�N�(h��L Ε�Ó3F��k�]�[)H}���0󍳡��6jԈQ­����?9��DQ�5��O5�P_��l+��cU�G�%��!���g�f�L��C�>zilѰh
z�*?Y�X2e#A�v\h_i�7{{*��ʧ�G�%��cg���he���蠘�5&�H���د��6~y�,\v�$W]���� %�9���m7�dZ�LD<L�Ur��B ���
���1MM9�<#G\�k��G���B�CFŌ��NľS�>EH�d5�I0˙Zպ��&"i8���J0���~P)��dg�
g�lJ8�tp�;՝��è��l��j|1s�I_����d�(o=�e��;�+��E�	�
�X������au|F�3�{��K��z�)�	���G�#��`@��j(��t�fw�m�I^�3\�Pl��%D:@-�G�r?o�喿��:T�rp��Ό�_���U[��'�k�����|�U�heV�Jo�?�9H�F�������4L6�\���"Mh�b`pp�j�1�kX~�{�.1'A<�;)M����l
���퓤0��Ɋ�͆�(o���8�n��t��Y�&=�M/�gcF���x0��/����1������;�;Li�����XP��ig��K�͸��n�����g{Gw�L��R�|}��:��.! 5��l�+��z�M��L>8����.xP?/��Ҙ�j�w�ַ���a� �,��7�LFW�ȉsϻ86^w�B,BI��B�!��#cΒ�u�3���TZu�N��jFrB�U��[�j������������ϸ��
E�z1�p����H��>?ţ�qjK9�1b����נ�8����(�cζ_�����G�-� ��,՝�pk��wq�Ga��, `8�kKp�X���##�Ր���\\'@���5�4��ofw�g�c�Ra���G�TU���������cT��"�N�_K����5�Jaa��>���&fAL��!'H�Ɍ��76�����U�ܒ�%5� Ö�����}�!��R�|�����˰n(	��oU��ɾ��q)ׯ=���r��OQy��d�I��R��� @�+AOL���L `=��d�t����؊�:�q6WфR�����2����t��͏�v���]��8ؒ�ɛ��~!�B�������h9�>L���ƅ��V���)H ���#iw�������䱚�x�:�!�s7�iԦS6F��a�]8!���Ɗ�J*�k�#��0,����if�6M�G��M�!m�x��orz�K���d��O�(+g�V|�'lf"�S�1���YN�G�n5.��AI1ix�Z���<f&���<4f(��)�'��pS��;0��&���A~x���D�~-�F�饿	�#Uw	@������]*��q�~�!��w�����H�&g���PKl�P%~�Ihn��>������i^��UoQ]2�G���%{(v��W���b���0���ݟod�y��Ѫ%�$u��=�
C*�IG�;�SRa8%�������,>��8~�fʙg�`��=��q�ʏ�T��@���/�`u�xꋿ��A([t�����s� u��۞�R�&�B�N��S00d�|�<֓������4���3��,�[�ͳu�Y���!�"I߰�i����Pw=6������뜖$�:�__�i��\�)g{�&�G�s���"�Sӗ�҃���� ;��T�n;>��#���G^m�݌eH��ѭ���!�6?���J���[`��'���΋>��0��2@�w,��
�j�w���UA�J�d��@�Ab�Gz^/X��p{aRJH/B]��2�>3�]�	����y+¤t�F�a���h��{�BsN4�Δ�"chG�^DW�Qj�椲�u�ɤ���]�^ע+�A=���C��	�f;�|��������j�iߡH'�LO.�%�P3 ��/��������Ta��;C9���@	��`�5ҹ�33��z��4Kx���cGֻ�AW!B��w������~5��5�>�7L�X�LO��g��?_|�Ր&�{�?�:L�xT �jc�iIϽhĹ8�@���$)b��MG	[�
歂� �Gct������Lt"D��b����t�h�=�$�2�72�"���)��7��9%��J�Ѣ�3 �o�;��U�8Z���n�
��h�����^��$�b��Q�g�)��yp��}iD��22!� '�r-s����*Kst�B���&�3���K�}a����$���N�EC�/�ݮ�KI�9�#����J��Jx-G4j��L��9�s,WV�����L�V�g��<,�ϲ�)�)ub�u
.L~�����f^��W�:?5�C�6/�<����},� [�3_�@y��-mo�����:>�$��`2��q��QC�Z����H�@���A4��Ԣ��V�$��E����zR�q|rZ���ܕ6���6��4�>�^��밗Ȓ�d�3��셖nBEI���̅�O��L��H��ͅ%Ce̎@l�&��*?�\�5dC����3hn&��;��P:�&�wꗱK �"�~˘�ߣү}UQ75�@Z�SЩ����D1W��]�b;>J��V���!��M\X_��y�r�~��7
:��0o~�!������-T-l�&��JK����p �{\�cp*�9�7����%S�m|�<��T+�5%q�z�Sk�U_�c#������l�0�1���l�s{Sn��m�1�L T>��$�Ә���t��;�ʣf�KSM��)*p6�$Q���g����`[�&?��������(�Z���j�b�O�9xȮA�~�ߵ��3�Gh�8o�r�/�G�bX�kwx��PN�Z����`�6��&�1��b�ee}� s7�)�Zf�O�Q�
�L�	��n/���˩�8�&4~:@�HMͶ~�d�ٞ��˨<���y^'h�
�����{�J�N�3@"n�B+�����,��`�RX��ǂ�[���]��[wƂ�p#����-%jA$v ���=�s0���һ8�!܃|�/7����S]]q(�-v�?9�Κ�Q��[_�Z�0:|��2�4g�����(�ߧ�2llU�Ŧ��w-�0|v��
��Uv5��I*�?�*[�⫑��m[��^��$BưacI��ؔ��$�h�ߤ6囋è�A�:EȖ�_I��d�t0��K:�.t�5�c�t~�}�.bC@�.txB�O�/��;W���U%dN�S�*)��	­ғ#;��EW[�x5��ve��,�@��dԉ�v�S��8��!՛D-�x6�����BM��Y~1X*:� o��&GJ�q���k?
a�������������%"��jV���?��>�u&�,�_&���.�G�$5�-�剽ۂ��47�뢢�����bxJ_����>�s�Ĝ+ۂs�F�;Б5C�&C���W���˄w���@���� @9�}儅�S:��)6NO�U�yN��o	R��n��D�����n�\�&�@�|_��^n�����Ce�a�)t��8(�9!^��'��mw{z)��I�;�Q�fs]6���������8�֚`A%4���rޕ���][a9;5�	�]��7u$�LE�@ww���U�30�� q��RR,�8Xg�!�[�F]�Z�9~u� 3ͽ�t�V���P���e~7_���|7e�u]6�A<6�NZTmi�+�'�0pz>N0Bs��f�T'�4T���o���R��.��0��˔«?}��C��VCbn��#S���5y|�J4	։���n�!��d��� ���h����k�r,�"}���F��m9��9�������o86卽~v�=S�ޑI����.���;�b�5��2{�m��=jVF Z��L�"-��r���(�+�*�"��:��e��K>�z!���&��q�J�����lS aY�* �@��)�#-���A,v��0��hc��z/A�n89��yl?�����a��	�h�,Q�f���nk&���h���d�Z=���<'r�j�v�����a�	�jh|�T�q��a����Ss�oeχ�FQpM	 M=��%��U�=��� �T`p�%�����G˓o��m��s���])�����e�0�y�ݢ�S�s	���ۺ�-s���u
�tpap���b)Y�S���J�j�`Q�G^1���ٮ��W*�g�ij=�3�@�[K-9��;���m5���:Zٕ��=y/|iH�*$��M�b��״� ��mv:���'�m}d�R�� �c�빫�CR;��Gw�<���T���fi�����s5>�,*�3���ug|c3�����U��-�r_J�#0�K��B����L��<��Z���N�8L��&A����or3b@?��֣wF��k�KBF�d#���;�?xO;zF���7>�=�8�^���%�T���n��ő|4-��2� ���U���*�tj5~!��#H=c�$-/�Ġ���m�L�-�'�C��-6A�O��k�}�ouh>���J�k��Eذ��ݯ� 2�K2�ϳ����Qhv����'w�D7�m�?�?�Ծlar{�PO�m�ʶU���c^�E�Sk�/^j#��kz�a�Ʀ�AȀ�G�5�JQ=X���y�yd���Zk��+�R��� 9;(	_�}��^�9��<���������}k��E����/Q�@zi��"�Fw�J���ώ��)C{��m�o�ُ�ǹ+WF�e�cY��t1W�r�z	y<O��B'vX�!qM�f㠫V{R��t\��(�n&������Gs��RUn����̕�A]�'�?�rН��Ώ̺(�^�~ǅ,�C�'�[�"L�چ��^%"r��泮=KӣD�� H�B��}M�`oEK����'��d��S\|+/�%�� �uit�Z�x#��K��T�w��!F�u��7�bEǐ�	��Ҷ�	�ʎ�k)I�u��V���)����������4˻��Kx;P��2�!�8�,���F�T*7�{%����Y�'&I�&'|��,t@D�^]S��r�58�{���R"��������-ݎO~S{-`����۬����@DEn��+��z���@��]h̦�@�-�jU'i2_)@�=.-����?�� <��	�X[
ux�F<�>�`A�tJ�����R�/|0�C�-��V*�d��W�K����U��M)� ��a����o��=H|���;L٬�Dz�E|Ļ"G����ݜ����ǁ����HhQ撾�P�-�P++��u��*���j)Ж�8D�H�ȷ�lf������w_�HP��=�|8�����U}�n��
���_.}���I-�^;|����� x?9�������6JB����8��3d�dzD���R�p�Q���q���u�@��M�P���)�m�������w �Ff�RO�2�eL�y��ؽ�¤ ����y�+��B�E��7���^�����(	5�G��6��S������ �z���x=�/b��׹ϗ|5��i�t?Ʋ)��D��K���C|������.�,k&��j6k��3`KdU�Р� $h�6s�~�[�'C��`����gqO�!8�0�y?DX��A;���Y�:�	�eӨF���7ԸT$�1̮���@�5o赛�4]k�i󴵦%���yJ�3�췶�P>U�6Ex�4�<��KCd֗�.�sy��y@��m0�h���ArX���d���8��� �Ĝ#L �������9�>)f-wu�5�t�)��N���嵓�DU�h�`}֘%�-��p�i)	��p�p�o�#5h�=۪��X�5�{
CM���ӯ��Z8���|*�'�Ipmw� �S3v�i^t��_�@������0Nz)�$�����R�~��6��E��社J�Z�Z^���P�+Z�4(;.�W���������H�t�T�K�#��B�S�ם1~>S��(��q�Yl�>����Y�<-:(P9�/�I���ls���~I5�@I!2��R����q�Y��#Y�9[^8r��:m<5?��S�/�ZJ�=�\WS�^����kQ����.�~J��V"ؼ���2��J ڔ���6DаI�hzy�{��R4�#�L����П���,W}D��*d���F�b�H\K���!��Z2��?��ͧ����+Z��a�ޏ�z���)m +��w��-礰�]�|��:%�O���<��e�0{zHo���<νH��GNh���&�/��rYƐ��erQ_�!=Җ;�D��^׏�[b3u�L�i��7;�;-\�=�-HV�s�A��Dr��B�[?o���&y��b�
Ʈ��ۦ���V^�`N�Íj�|���2g$ֶ�U���׆�����g7x{� z�rSA��q�$\�*�ӛ�g��Y�f���A����w���)bR���zT�?@�<j����$xq�uS:��<�v��0,�:��:x&z�2r������HN�+_���5�_ ��n<��-_��]m%�����q�����)����=�DAށ�R�N	4����\z@�6d�9�t
)L"��.<��d�ެVƊ�=����=*��Ҫ'�:3J��H�{�[l���T ���PJm����G@������&��Ν��pb�O�ÔM1��͢�b�/�����h	���Jn�.�P��*�4��E�����H�r���A�p�w�* .��E��EZ�/���+�ʆ.�x9�K�>���5d����?�7e1�.�ԥ_坩��{���4՛�v6`}�D�΄h/-d����)iu�m����qp�g4�2c��rn�zٓ/����2&���$q�foƂ�I[60=��)aMU�r/���ɲ�?/��N�5;[Q乙;8$c+�S�����Oخ@���^/F��~���<?eᡚ���{b�h^i�Y�� -Y�8��OZ��I�"y#*�N��ȑ�v2�>����ӭX�� ��"w�1IY�06���Y����[��tJ)C����7輤�2ҞYQ���w�nUK��[.�ﻡ}���=��Xd�-Բ�0-�J@E�ݑ�6Sh�u힏�J��j�h��z{֣�7�4x[����A�ץA�=̑
���R���l��=Ӌt��j�3-?Hi���"�lZ?5�B5��^�"4�Ԇ�n�Lj����W�|����!Z$z��C�#>��j���$�v��A4��K3�S#�wU�{͟y����sx]���x�Xs�s_5{M
����͐�W��$�<��
M�41�d�U�&�X�� ����HI�s�廑(�2m��q�����ަ�Ɔ�Ií�Cr�J,�Zq��Z&[b�W&��@�qۊ�L3�WcS>��.�� �5����=���Z���k:�뵪^se���~
�5�5���8�N¥��h縝Z9�:t�r���QK�f��@��2<�z���,J�i���L7w�c\@�7���%� 7$R���cͤp/N���\�{kb��l���=bp�̮fN��@s*2JތF=W2�Iԧ�\B>G'R$&��$��<������A���r�6�Td�XL<ڷ���ް�U���P,Y ����!���'�R�q�a6��dP3OT� F��"�B"JCc�*3ޠ�L������n.]cc��"
T�p���,�)��4���=Y0��\��j�n���b���}>�a �<�4�ʀ,2����Ժ�E�3��
����f kS� )H�%=	}V��f��yM%���l��0'ѐ'���bQ_ц1�'���vk�h��f]KOӑö�·|jj^dO�x�9�)��Eu�[�*6ڝ�����OH�A���Ǔ(qG��cZ9�έ�GmE<�hGhτ!�W+4̏ ����%|23A��}'�XA?ү�`��i&JN�y�fζ�p��	
�'�ގ�rj��KSC���\�9�[���v�M��{$�e�XX����[��c} zţf����[�m)Y��o�}�@FB�+0�������ۼ�������㿗�J
+
/P�;�I2&)>��,�L� �න�"A �۬�3�4��?�W9֌\F�������:��16�y�f<?^�;��߹=4r�h�Rf����c3��g����<L!�zC����"�+ߠN�K�PG��[	h�f}9VsH���CcC2��ހ�-|*N+-�}�w.B��Wf�5W�;��=+��p:�d���HX�^�/��D�kp����7�A�v6y�N4M�#���O!�=��`��ʼ"3����l��{Z���kƚ�uyq�i��I���.��[�B�wz ��,]���*fhY���.�T��.$r�H�rt_	�0�۞������}�W`�R�27�8B�$���2�3n�OU��M}����#<�ycK&?OR}��-ꦈPfV��AϦX��/�����PHys��.t��a�%���E��Bp��#]���	G90��b �q���%���o��l ��C����G%�sS6�$㏨� �uxc>�jYo-��!aFj#۲�y/�o����uM�����.+E�꤬�� ���N3�B�z���u.���k���ҹ����O1�^]�H��K�'�3F�����=X��J�}P�-�P��S�	*��C<-��T�Vt�(�=��
��?�|Oٌ5 Ҙ���< 3���P�hu��q�ז��ϋ�eGsV�·)��p���UT�f;�D��n��)�����&,oKl.g���JyS���/���Ĵ:��1�vv�撈7'R�Ͽ���j(��cN#��K�2�2ꈆC�X����⹯�:��oʁ�2v��;��i<��+ ��y�����QVbKOe�R���V��"Xk��^Ѷk�Z�ܼj�R����XfF�a�K�����A}�M��u�b���:3��M�3���mheE�I����Ƨb!u�fռ���]B�>8�V��s���ڐHꇿ�X0�����2��j2z۬;�pG�6�5 A��X���'�n&���X5�M )ǀ
��j�N�|��&n9Ե�,���m�N�1����KK)���>�J�0��!� ����D�d��h�J	ڶw���Lc\<�;b3q�d�H2"�Q�BI�c$�щÒ^���J
r� �{JG��1.���\̞l�)�8�Eɠ��0�]r�~�e���ps��/�$%��T���eoS3��V|N�w.�W���������V)�����dw�����L�@z4/��>6my��޾Q.�M��S��)<f��7����KrB�;��a�� j���	g�o揨z��n��O�V�V��.�B��*�K�u���7ġ��މ�^u&gb�A���j��xU�Y�(|�E1�yI*�N�\��q�n�H�2$�1�8l��}��L����FQYN�fx���/C_sR������V! i���0�.�/����QDi�G����X��RW��_��]-�0�x��t��}8���*�I��H|�{��+��24�
c���8�'��cʒ�P6�fߗ�ϩ�'￷��k^�~�������yÛVG�4�$p7���[/����?�N�.��9�R�v�&;J�0�Zp��%�'x�s/���@�Dq�O*9i2��"~��Ѹ�F��v�	�����ş!���@�G"��>(���p t[N�i a�}n92ѠDR�N�d�8���!Q�OX�;���NZ2��7�f���\��Ϣd�Gw';q.viN%S=|�v7��c�u�UIT�0�{Hz��|�x%?�H��]�Oꦥ�z��30���aR��#�6T]SZ; mCg��4kax���y�l����9=��RlV���<��d	�Z\����p��d���������6V|����$�& �>f����R�#^C��ܡ�,eX���w���GU���Cq̋��%�２�5��n���H�?��r>����C�)H�q(iQ_�φ��@,_H���My��<U�X��KU�(!�+p���3�4���=�L���fV!#��X|�]�h�)a�
i���3kl@�������FT>A�����a&G8�y���ւ=���	����%A���M��"�T��iy��͛�3)��v�K�M�p"O��9��;���?��&.��&j�B�n�[���9*~s�s��>=�
�k9����Z�8]
	�uP���y*-@�����K�YRC#�vw�Gw�/��Lee�ٙCY��G�`lp(��������+�T���{���)�x��9��6�V�ҡ��ěX�C����X��ث�/lɃ�/k���}4!l�I�V���)����s�k�ՠn���Y�3�s����E/Œʰ�g�Ԫ��Y�&N���-]�@xN��_�E�
S:=��Iq��]}����R�UXܸ�I��I�"��Q�D���L�n�fѵW�1����\w���T��`�{�
e���@\v�r�5p��Z=�^���ѩ���VB5t64;R�P�K���XI��8-�h�95ʈ�����1��8?)S�O�؀i�S��#!�4 U�:�ET(=i�S]K� C0@��o�
�i���C���A���\���3��|�@c�X��҉��Q�F��&��ݵ!�Q�c��p�+�A(��ї��V&�T�{5�	Z��R�J�#��빃�uG���SCѴK?��wYF�}سP0h�<ŭ2-]N	s�mS�Ssfy�!�"�1��g��Z�ᢚ�iqe�fN���\��a0�e��d�����6j����Ц]������{�:��R�P}�<�_B �~'tL�>Q�Ӊ�h�f��X�q��Ι�E�@��k��$����7�L҄��9� Y�@CL��L���h���m�p��~09�5�1٢���{���zL�aj&d�N�L``����,(��М28俑�YuO��5��-`���齕�Q-��a���^�������n���*,�6f���[7� A���'�,5��� �)�?��&�W�Z�>����D�Q�M�d���>����еh����g��׀k�ԹE�,��d�xIpdɔ����M��ov0�;�ن,@K���u�40�^�����a<��E�\7�O�3�g���O0Z�@���0h
�EoL.;͝t"�Cz������fR)��i�?|�.�����s<�b�2;x�������0/�X/���G?~9]c��w��m��@l��ƞޖ$�<�7�>�gcx���m|n7�8�fF��Y����Z`����e����fxE~j|f\�ѻZ��l
�i/��?�Cd��+��1�Bv�Q����RU�eR��s��J7���I�L��?k��uuXw7=r3'�1 �SiO����9��8�pŞ��'P	���%�*t1��R���!!W�.������'�␵��+�PG9W��:BR�Sk���Zv:���W/����� b�@��V������L  �W��"���Q«�܉.���"e�%�*h��rל,���_�E�_/V����7m�0d��r:J�Ly��msc��ux�֚�+��L�L�JF'�b�+?�g5�+%}d�~qCz~ˏ��ҿQ;%��5�}�ڳrf,�@w���l�/����RxP�{����R˜2�%;W�9'=�� ���e�ĺ�s��v1D���b����%�%��1����¦Z@w!���l���_[����g�Z�p##0܇���[���-7o���D�=�s[u�Dى\j����b���d��ƿ�,V��
-���Gk�3���M]�V�M/=�d�mI4�H���6*��]�� !%^��5�vx�$z|@vJĔ�1;s�J����ݖ�# m���v)��K�MQ�*m����(�N��I��!����v���n���PR80�g�{T���Ҁ�n��xa[��X\�A�Z`���&��;s��:�vR��ey��}ۯ��\�0Zw��쿽�$1��H���Z/Y�![��#dF
��Kd������`C��/e#i�#����+j~���g8�N�ך�O~{����`�ݝǩ�@��H�X�� m��a�v�;ac����s����gh�����(�N2�bƺ��P�8s� -�C�w�-�E�4�I���ϒ��}p���N��丟'm�K��),��Ɗ�y��`���BҦ%NChZ.���k"�Wt�g�U��|�5|�c%�c�<S�I�B��h]@#���m��LheY��e�� ꦐ�v_&��WjLk�FX�Գ}��NZ���ϐ/gg+"�������/�]��U��;�����_��_��-��C@J��М.y}A����j��k0�����#���p{��6�W+��C���Q킓��k�"��}�z��*B���*lJ����忀��w�
��-gL#�xȤ�1+-)>DQ4+4�.Oe(ց�J 2c�,�t'T�����]�`���y��/KV>�`���[%폢'�]#^auU3�D_�3@��/�S�x�M�{�g��'/���x�����h�F�#B, ��~�ڦZx���CҐV���b�*ǜ�����c��Z�~��߰�d�� .��`E���]��]���bA��Z�ƍf��%��^A�%J�f�g�F�˲�:
5����ǀ\��T ���+e{ŰF�\�ukz�d�[�"�dS��N�+�g����&��K�Y�}`j�a��8A}d�X쉌��QCmɃ������p�����d��a;�	��u���`�~L�r�kŵ(�+�m�؈g"�ZVvqY�0�*
j|�V�8�[���!���*I;X��!��9�y����̟�?1��r�\�Q��9�5���?r���?��F�R���[���q�|p@fl�oF��c$0�h5���N��fD���8!"]�˟����e�����=�m��S%Y��2��(�Eϊ)�Rp�����_0i� ���'X�fE���}�PLB�\�w�^@�6�#�l�0�q9�Ss���`·�YJ׎ө��S��S0��ui�����Ep�ƍl�Z���5R��!�aQ*oU�X�7	)���DV�ie����֥���e@�8����{���� ����꟯Il���КZ��>�@v��󞐲ߛ���v�%à6ݠ�4�=%^NTPT�ط���/q�ߡ%w���Fn��t���T�Um���9:J�t�g�yx'�4�ԝ���H��7{�ߤ���w+GY�
�>�,]6XO���L�5t�Ms�����h˪}�xo|��(��|�N���Ne�8)�i�1���e�;��ӛiۓb���v���24w�u��~]��.�r�qN�X&�Cn?Uz��(�X�e,�T��;'� �}�Rz��'�=֙�O?��ja�#�ȭb�"��0��m�jÇ����>(�����"<�qws��Z��B��gl;%�'��#�,�Љ����{-��+����f�����"�.O<�	�I��X�W�L�@!��5i���+A��-8����M�@O/�l�:c, �y�Y݉J�=��ׅ@���f_Tߙ��$�xi�r$��]��M/K�*s���=W`��� |FX��͸�:j�84.��}
y	O��ty����,�`NU��~�4�<���J��h�=�s�A����A�Q7��c���nN���+5����I屝�¿1XZF^��g�`ې�hk:���� -t$lt3�	��=,�9��֬��H�H��ztл3�6et5��f장�8��d��#��h���G�&ASy�D6�x�>�Hk����N�b��- ˫ }���O�����QyFf��*�[�Vui�xV=r3`u����oTdݾ�A�n�Qm����c蔠�C�#�3�H��せ9H��򈰵Nmg`P�䊈(�e���Z6�#��UCZ�)�ԩ���K���/������6�j�s�ۤ��C�Aͺ��,e����d�P�uN���A�L1�w�i_$͖�,��輅�\�
\|>�i��B!��U9M=$M�9)�"�O��E�ۿ�8h/��(d������F)�>��Y���ͱ��<�%��\��6��}��3��c�|'���8�:�>�gD����P��E���*�#q��r�c bu��~@�J�%_���FIh#����=��V�%���ϴ��D�z��;�+�`�;v�8V��y
 ��4���.X���^��������<�@^d	G8����k6Q��S�%S>Ժ�-�޲M�ƙO��씈�������g���G�HP%��#�-E��:W�U!����4�7�0��ȼ�a)�6�� �ۻ���A�֑�,`�ZͫP9�DN�t��	����z�4I~�^�"�%��G"t��]�<�Ǯ�s��� F[x���`AE�����)�T܇D�>�Ћs��ȩaX��W�pF�3�d�r�p
��;����(�Y�+���1�1E��s�>2��!�p�ۗ�����҂����_ �N~�VQ�>����vAC-f�.�Sc�����FE����񆲎0������N���ډ����w�h����BN���� O"�L�Λt*����O�i7�WV&F�!�Q�)+eq�SZ��Z�U�͋�z�fᎡq���'�Q�~cTrnC�Uw��k��3\�[��N��,��֮A7�$6+��v������[e���2��f�g��C�^��9���W�,�V�x�q�$��n�eq�7x9����u_$	���n��(�q@jISv2i:�;�k�$c9[hI	����V�֓��*vg�|����8�Q4)5ŵa������|����r.�~����ϕ�
U�fm�q37�W���k���ڵ�%qA����E���y�ٸ��x��h2�	E�8��EzT�=eE���a,��+ӿc��e�4~��Ľ��'l�U�0 �QH��r:�S+��d��C�`�?f�����O%{�}W��4�Z�����I#wd����[�� rG�c��Sc���.�9)����B\k�@�p�>�5(��;GVvj��N�ҷ���]Z��[&�x�S`�����h�Td���1�Y�y
��',Э�sB��.m�E+)�0M�c�5�v����6�Y�8aC�5��Is�+��u%Z@�7�ǩu�+�����t�W 	�� �+�T~^�P���;��4l��=�K���%J�N�q�����	�nv6<Z��9a�}�e�I���U~��.jV#�����?�|�����uy�.��T�Q�}�:��+����밈_'�{ƈ�[sky� ���dP�X�q�XLۘ|�9����G�ʵ��s�l:�]���`$���J��/�Q*W�*�1�o��nI��1�H�v���L�us�ڶ!}�sf���j9�Yj �.�>ae�u���{T�ЦÆl+��>7���w~̓/P�f]�ˣ�|6��YDK�W�g��Qg�MI� tȗô,y�#��|~W4O�K����/��nL�";b��2��DEz3�n���;��]㮖 �2����)O��+)���"�þ܎1� �]`.��~�E��/H�(Q:1�s҉�=,xM=<=/�����)+@�I!�I�8�8`�Q�p�4�&$
����q]����
���_KN�+4��s37ʑ���$E�Ae!g���_���y���b��=�v��-��)s�C�,>�py�}��yT�[�~�?���'����XPoB�KZ�En����@wR���W�GX�Q�O�=lƄ%��S��U>�~W�,sk�}:�"UG�Y�<����n�9��I^N{�CƹT@�E����<+O��~NL|[Y�dd}�k��M�$�����B�G}��Pax}�D(-�7�kC����ϲq���Ҭ��S�c�{�RZw�h��Gg��1���Y
7��3�<�F[R�;�m�Kɯ�=�����")��צ.�|�N�8)hR�A�6�s"	��l�c0:#53�Z��ݙ����ۤ9���������mck�a�4w7���s�X�F����(�M�S*��y�sۢ�\1�X��cev+����I�����y���GF��J�DK�Ӻe��`#`�Le����U$/���,�'⇿�P������W��n�B�̹pKh�Ϭ��:da�p!�t7�ԗ�;��'��'GW�C<[Z�CV�{�-䎤���}M[�m\�[2|����\��
���S��°^ޒ~���k�����4S]�ع�ab��>�V�y��٭��sj���~�hU��+���6f��?�.� wHH�0��>ݰ�����
�N0�܇�sۻE�	N)����/}�&qrܢ�VB�g8-�BV�J�'�2�c���i+��s����;f�b�geoU��)I�]�.Q�����85~C����7�%��5N�`&��U�O�HRz�ٍ�Vӕ�a��>��p���ҰC��a��K�}�l�ڤ�H1����]�u
޾���������J���&`�:AXM)��X�
Wpm�2�
�7l9��$�����b�ij���O3`1`�Hc�݅ ����p'�ƺ��RWn�<��О��e;��@�He:*�DAK���� ��"�f+D%I��
�eG��\Dq�����~2�C0}�������t�w]l��Gm=B��|���P���=��P�P}���M�tw�*���@�S0eۉ>�F�!B�{���X)���3dW ��>�9��y�_��/B�B:�������#��>�����j�O�T.�0�V���t�����R�H�f�^�Zo��şgVCQ������:�W�nMWH�󲭿𗕪�`����	�d�f���!��G����e�E��S�2>A$���XOC���z~I����[� ���e�4�y��F$GmIX�Zѩ"A!C��6���v���,5�|�3�A��s��Y�N��n���S)�o=#���&`EE��/��/��Xc�]�}�����K�����y!\4��ʊ�8��Eѵ��x���O� ?)RmNq~A��,~5�1���n,"���?����u����o"x����X����1�˛�㝆=�}��.���22
u�W7�a5}hۨ�̰XIDB�B5,�9�	Ӷ5���E�i:��	�-�>�m��[�ᙘ��[~ m�aJ��;�b�p�ېm���J���l�aq��b�~��PDC��e�������^qt��[w�>ܿ��a�4��ѷ�/w���`Z�[Hͩ�T��=ӏu"����p�L"�)��8�:�7(��)�F�"Am��c�عj��8Ys��d�3Zv�H�mgk�Z�<��nr�Q`��-gk����'W6�t��LK��N�q��a�7���j,s�0���c�F�[0'�1z�c[��*Gv�X���� x�d��Ul}����'�@s�!�K��4�m�1�$��ې>��$�ƺ�a�_:}S��L>���GV�C�[R����B��a��1k���-z�h\�Z*=����ל�2�
�w�¯���>��ye�J%򳁷��_��D׀ˬ���H
�.�;*�����Ýc�t�Q�aoM):;w (��Y����8��Yhu����֗�~祬���;}u��@kI˨��ᲒdY��?{��%od~ӌޖG�?F��ՃZ���+�5��!��G���y��3�k����TM�Y�����{w���h1m�\k��+����p4r򂛛r�`����)u�?�0�KP�e�Զ�f�	���(��<C�#syz�_�;�vp�x��BC�U��c��1������3����<��&�k;���%������տZ��B=թ���C����\�g�!���by��ol���
F�w�� +l������;���'a�R���Y�ʷ!&aYH�3��}��K�5��'�a�L��v*ש�=:���S�ShS`"��,��|W_LW@6�J����ks����!�7Y�?䥘�'�R  f��&[q=��Q&Ĥ����&H�V�l��^j@WNa���ehFv��i d��5TdE(?S��OO>������-�����y����:��N�۝���{�Hic�^yǚ���v���>��&G4�\ ~\�zp��8W�G����<0-��vs�ϭ��΄x�pK&-�4c��W���2K=	�K�R�3G�=/�0��Z�og��3���+ϩ����-\a�޳�{Dái�۹F6P�;G5���3����\���H@�K��\ �Դ�˾�]tD/���bL�cjx���]B�"5u�̢_i6��Z �};����dl<�L��%�>F��ib�o��cO�5F��e�sWM<�����@0Kô0���_�1F�{-ݨ	7
�v�|��ĳ��pS��ܩ�����*֊;еf�1��߽f�x�8(͎����'��AF�S�V�yT��|�j\�&Q��n����[�26��j�PmBB (�֫����+�B��ӂV�K�����h7ܼ�ͯl�pԩ(�oW�C��m;�MX�dL��� g�c=�N�������t`\nۿ0�~G�}�,`��J%�����{��&�F~#(�x~G`?�~
;w�fT7�t��Ǆ�\9���p`�VLб�8������pVG�ofϭ�P^��]R�L��G�U��V$���Rk�Gc��ʩ�]��?,YN��@3H@�Ţ-�[�)�ļM�����Z�0W���zd��mǔ�GP�W���s4&0Q!�x��������g����ľ�Z�kGK9:D�0��Rۙ�Y�O�0lMh%9Xyn���H��E�j�J�EzE�t�KK>� ���lF��Uj���öm�/V`��;�jO׹˲�3D�ET�V����Yk�sB�YOF+��u�%;�=E�VO��+�^�U��g7�l~mwV�M�.���V8X`�������_��E �1;��H������F��������[e����)O�p�p(�0SWr�GWM[ƥ��,
�Z~g�m;�y���wU+G�( �ڰUI͆-!��6��k�Г�~���Vs5eEﵓ�����v׉>C��Y�f�X�j7���˵�,U��E�V	�������|f/+ɇ�,p{k�=c��"�:9�EJ �ݮ��9�{���Қ�����qa��u\�a4�Jmg
3.��A��Q�%�x߈_�ϊ%#�U/�sc��>;t�8��y�3G�?\`R��)�}Q���5�=����(�~P`�]���q-wKQ	5yt��J��`*��u
��5������ �/��we��_�J�\&��Y�M����(�L5<�ƛ�3_p
����89R)%G����P�q�}6�@����4��g�c�y	\*��S���x�2�"���,�׾�����|�h�G������'���C͝�"b�P�o�J�� ]9�������a�Z�p��j��Gr��^^��vtD�&u`2���OAz}�`���%CpJ��Ps�>��<�b��E=��]�'��T~�@��'ݬ��#V�f�n�[�,>kl��x�߱=��Z]�G�,���?xʉB/%oMǜ�!������ghW*|���e��=5�o$&o��f��JR�"&4.tx��tΡ�-G�Ks��R��R��L�v�[�EC"9�}=� w��c�������v։�:oA�r� �I����������ȸ�}̹Nz4���JMN�dB��?�n�ft�����'v"}zɅg�/��s�O�?��+���o�^biVP�������K�1xB����p$8�W�8 A�֬��wE��c����|��o�|#<����Jp?bv�4J+�i����q�)ç��B�
��}e�iu��Ɨ׈"�Fn��3S��b�e��oH�0%�q��í�m0����G఻`���{|U'ξ;����J�o�S��^�rx�(EC܌�c���p�A����]Y�=5j��5<Y�4�I��b���%���"8�T�T��̬K��˲v���R	��E��M?
|d�)���\���Aƺ�+����&������JI��62ɶþW���'_�Z��eR��W�M�׏'����~��ȭ�8��~T��/��-��O�N�@��yE�a�mE�.��ҺVwxoi�b;�=�?H����N�f+p�ۂ�#g�,L ��B|�\E0�>��Ҋ�/
��,n(��C?v��"�/{���^J
��l9���V3p��s�����,(��X{/���w��� Cp�L��-Y�.���	����'��ج`}���n�!�R����~��l з�I��R���8h�������,ϵ���fj�(z(�'-�+�1��(����6���ɀy>�;W4AI�\��nO&A���&=�:B�R@$�&<̭�9p���kݣdR�9#?�]��BXN۫�d̄�ƍH2p򗘪���I+E3���W(a�Y�"h���ŉ��s�����VY�����ӎ��*���iaһ���,ot�6}��qCg~��d+x�^���k~La�_�4�9���u�?#�����>cNnU�O�Z�ur���(�7
42�4��aa��,���A�G�OO��c�p6K�ˈ�d3%9�������կ�qN����z�FSK�Hy0��N��s�T��H��r'����$�a��PkN_?'�Ǟ_��t�^���8&��)\x}��S��Xdi�������h�ݺRH�_��eI��T�Ym|���c����˰
lN���CW���k�`�!IcԎ�{�8�δ:N+7o�LGHdj�`�*�U�y���&���{F���ǋ�>)\4�\�9˥��' �B],���,�4�w�
���͹��fV�&:����	�iu߬�	�����#��;���]��Rʣk�u��*w��6P����7Nb:�M<�/��^��B�hE6��N�F����[�&��a�^#�W�>M.��~�]��~cv*(k�eZl+&�b��-|��+��>��������ʠp��e�a8j�UЕ̖h��Ҟ��3}�5N���4���/�a��xa�5�L2|C/M�^�p�_�X�	�Kq�.cx8u�e4:cţP;�.�Ü�{3��&W[n��Ԓqe�:�Nz:_�<3���%��`�ə��8)�f�y����k��f*0���7�?�Z�1���(p�l �ͺ�c�*5���#\�dt������K׬��4�
I�;a�T	��T1
�jj#��|�����k�>x��l�}�JM�Ja/^����(��D�G��.>�'�m��X�	�ǃ��S�w�(OO��[nT�Q�ֺE����:OI\K/�,@�1����v������V����/ (m���Jf	kغ�z%��E��do"�E�=ht��/�񛆃�c�9j��^����U�S��C�$��Ӝ3��O.��a:����^$Vȹt@
�-������*����z�qt-�JQ0��)h(UlA���b2o8����t6�'(���Վ>��c��>�����v�6Ek�%��AqW��\��H2Q�A���Hd.,�rЪ�0�!��x:����~;� ���r���ZcI����h�bL��J움vSb櫢�ԏc}#`�B�|Ei���C�]�͎K~���lZȺ�88�R��G-��SY��i�H��{�3� 1�6x6�a�%�+��㉻Њ�2`�>zǛw}���4>G��;`�ވC�� �� �5��@魋�B3��5Sc���a�c.�M����p����xʳ�m��Q�/4��+I(�!кT
�u�+iX�����pM��Ny49k�@���Om�ʉ��%��7~1D�yS��e��.��ײ�=ߕ���(Q�T������=�-H,��	'K"��
��3?���P�a*DsV�u&���#0㣑FR��9%c�
�-A�)�>t�ihg�C5�y��_���"5����ATQZ
s9]�F ��I�?�D�5���ѳ�/(z�z�h�	5oiT�q��pF�߷���X�DkKp�I���~9r�}�PCOu�;��y~��ZcͲ�z����G\t'p:	��{�l�!�%yk�aB��^�!���Z܈�P�+(����]�*Q��>2�a���d�nf�D������;q�p+��7)ں��ؑf�KQJ��h
��Hث�$�}�k���C�(��U�ÿ́d\���-�����CeB��J��@��o
�P��*�=0I~��o��6Ĳ�E�>�QAy"��}�Xn*-k?{M: �����1�g[�N�ug�$��Fl.�UV�]	[����>H�R3��(���˗'��(����0���P
�e��W��b}d�$!�z��C'���{y�����Qؾ�U�y<	�SD���I�?�ZzR�%o���w�1d#�U�}��)��v �t��.�B�.
чO��b�h~�;�6�{���Jwi%
ږRE(��t���Ж��רA�U�"冕��e�+��[]Yçx�-�6�Ǫzv�Ac�/B���t��F�ik�B�]�G�k���N��|��|�����S����:ځq���ݬ�׸�=d]\.�	��h�l	���y<��@S@X$`�NS���$���@��|�So�i�V����}���bb����C&�9���N�ۜ1������W��;��i�0�^~|:�f�KQ�F��@�q�+3�����N\s�=�|5��J�%,Pr���Ml�)&��J��(����"2�B�q�T43g��n��PS���vW�=/�����k'�G[c���qv��x9%�'].x�����}�䶊\C�]۬}�?"S���*S(n��ћ 4��lΜ�p��|���A�%㒨�P<�u��}�bYK�fXT�Zm������c>nt�Ϡ����-C�3+��p�N�B��s��:���N�\�v,�5���XK�<q�n�%��&���P�o2`���|B�L��{���2����A(z l_�0��P"B��ZMjd&�	]����>.dQW՗���qļ�v�_#I{K����_�^~^?�+a� V&�K<E
�O����ެ[ϧZ+U<���8�S��2�����6�6n-�I�#��]G4�O��w����D���gl�24N]{1Kļk���H�����Q����8�	�$O�Ӡ��ñ#����*�%���Q9����_�^fD�ml'���O�����2HJԓ }�75�Sa�O����l�?yع��5�*�YV�E�f�7�]�4�/~hq�e�b��F�('&b�K�������M0�j�o��;u.܍L�����e�ǠDp,���$2�Y���,��F���)(o ��)fM�陸��i���HC)���ִ�~�JAsl�(�mۧS�~�pK��2*�S�� U��
�4�CeQ�bJ�nϬLR鳜��}N��J)3@��]���Et;Ӭ�\���s���T�&�!�5���)r��޶Z}��E&�Z)[���*k�[v���q$��1MW�ؒ\�B�SkZ��Fj+�]��wݱߚ��\ޓ�a-Q����锵	P���{(�q{�(8������]r^F;��Z�x\�~[�"^�2=8�(-�t}�M�����ꨘ����>o��.?��P3�����kG�|��>֓5�]eQ�i`�y	�9Rf�+����i�<]��}Nm�?4b��rt%�jcBC������{��~��PO(zA�hsy��]m���'~��,}С�{�@�Gؚ�S.�v(�tʲ���7�����U������fN���d+8嫌=�sp+�)�	��*y>:�Tn�a��ɟ��_G�:�J��s.��YŊ�88��r"Ř
�=���9K�����u�1 th�bY)q��{5�VN!vF@�a;Ƶc�p�a���?�l���n� �������`���b��q�i7)1,�b|�f�A�,��m˦�7�^���f%�7N{���@}3-�lp9l�|W����c@�c�V,���$��o��<��_�o�z��0���Y�GiNF��&S=����$�/&�\�΍>ʚ��Q����+�C%��=��ͭ�-�d�T`�AZ��7ҳ�y���F�� �OXD��VXj�
��Q2f��r�Wƌr+v�9��FHtnX�y�� un(�C�����޻�6/���sD�c�g�z`�YN����zoP�U����yͰ�_ԇ+����x���.w������t����
3��+'k-:����!�R�o_G�Þ�zѓ`�������g��HGWY��՞��:BP�����b�ī+x?���	�	���]bL���FZ�Ή�!w`��.��Lㄳl)�ɼ ��j)�������9*���R�&I�Bb
+5!�iޒ�;V8 `c����rP���g�
9 ŀ,�J�<��ԍV�`p�����=%��JH��,}h�Q$��j�eTDN��0Y@8��hlC.�mBZ7P�5+�;��l����)�V���Ә�fIv�o2_��c�����Ɩ��@���P�Y�yt���J��:L��1��W '�H"����qEZ�q&0�C�!�K@�\���j��"W*�+��a^���ȫ���Y&^U�4X繯���q���N�C����[�M�8���{|��Uχ>A�������� m�����V�^8�N��ր�" KN��G��	��6��:�[^���B���f.o�k�B���۸.&��s!{��Sԙ����Q�)"���T)kK�*B�N����P����YY8�j�A"��������۠H�C��pd����5 6��% �!����R#@�;�TT�:������Eq�T�t�L���$�0﶑�8����v���_n�1�X�
��wq�
�!
j/cWv�в?B���~�0�[T�ZQ,yNڮ7���)�{C穩XG���|��V����d����nj��M�n �LD�~~��<����!��!|�А��p���m�ָ�n�?�X��0%��v���Ҩ
���}��X<�N�-��bh���g_֍ �	�����0��A�2�w�g�/�p���I�~��	L��3��S�
v�_�yH|���·�j�q����N$���m�p ����ӄ+�z^
K1o��(�X��0/
g
��W�p߈F�O�wv��j��e�Iu�*4�ч�T������D#ހ�ć	�k�"���+�L��K�������4����'�d^�s�ҍY�G�v��=a�����$�܉rPm�P��(��\���W�ŦQS�ެ{� Ymz�m^����l��Mݍt,꼈4Ǡ�;��J����4j|o�"y�\��y��Hy�Hs��Ó�	����s��O(��e��v� ���<ol�w#>v��5��KFI�c�5����Zeؿ�����=m�C�t�T�M���\�u�`	��?�B��{�C��6�%����p�Z�;@��X � �@ �b�|-���9�Q[��/��5�Q�[�9h���$��%0��,�ܝ �|���S-�m#�s1�C2٩�-����4#����ld��� ���FL���铽ݳg��,�r�sqJ�� �ڤA�q�Bz�"�wX��{VU�R�&��h�&��Yd|��r��p1$tYtF�|O�5ԵݽW�y�#�IK~'zY�USi������h�O�_MFnE=m��L�w"J,�?!���/`����3+��:�`�vK>��{.�D���l�(�CB��ɑ�q�M ��� �J^���Q���Tg�`������b'ڔ��}�r*��ð��.}��߾��/������E�����n�������2�{��Cx��e�g���H��?*ѡ��G�5���(�Kڣ��ߘ��r�8��}�-m�M'u�����ԄA��^�U�Y��ku���	2@���VyT��ܹ�BGL�r�n�HK�]}\+���{k��y7*5[Ǆ��OȲ~Ô��w ����=��u`��4�t�֒��~���ɟ捯4R���_&�� F� |�K�X���nT5�GR�
��M���p7�%�Jju��ο���� ��}�)�@�n�P��3�n���#)����.�w�a(�`�L�]t%��Os@�'RÊB��Z(�k;����-�~��S;����I_!O���4�Ͽ@.@꣯����7��E��&�?�UHx�^rI�8-���hV��	rA�x�5�S#�3w+r�����T�yP�k��jn�9����ab�!n�pL�M�0��~1���`�vVp�C%�޷D±��m��r���b<�ȢM�mA�z�ϼw�c瑻I_T0E�]�(��܎���*��)m�t�,`��}�H�o��{�)5���Y���}ϑ��(G��0�is���M>^Vyylp�<gj"ZP
XW�,U�;  ��[f�����L8�	!� �X�K=��P�*;���-c9�c	:�*f�ֆ�r�$	�?���H@'x�6�;�Q/�)�//x�\x�o��K/���� X�?9�-�3�tǤd���[ߣ'���Y�_�俾`0eF]%�o�@�]��r;�k�F2c��z�OgI�<�l3:f���8Z/�$Ln��ց�.�Ʋ��dj�Yw�ǘ�c1e�|^�	�@[DMD\]�bď�`�z�y��"��ϒm@5@�H�R�R!L���f,��dJ��șo�Xl�9ʙrީg�����.�C�Q'��׋��g���u��� ���̇��������(�4�K�����Q�m Pw��:���))����w0}6�J��Y����s�+�ԩ���8U�z��SE# Qɑ�Qw~�,�X{]�ٕ����&]��n�;�d4M�&�i���1�]KVz���������GP���mA�J��ԅ�Cȅ��LN��lx �Ibٟ�Yv�tx���G.;�]��;8�Ek����yQ��Z���;s/Ώ�xOn�|�<�#�ob7vb�#�l`ߓʪ&��1�G�\��#3�PV8W/S֘�V|< %sM�͚d+���w���Fy��|�֎�y�~�B��`�D/���򛷢�3�ۤ�ο�,�(d�1�?Ѵ� �9�$��B�}Sjx�Y@p���0��R
�E�ܩ��dW�8u*g���EϜ��& �7���y�#$~��"��Շ��T�TF�˯��{��z�D�b�b�'�*���d{k����3m�^{ŗ����_@�>3vp(8�Gr5'���}�|���C����|_�5�9"�{���=f(��|"�U�ճ��9�`�qG>�w'ܩ��R�z0�"��]��W? ��Z�(�h\ϸN���[Һ02�[o��W���=�?��̺����	�~e
���������{B~��΢�fn%�V�C�>1R53��E��4կ� $T��׷3��vx�X}1���l���%�/ym4n�z��^�u�2i1).��~�ԧ%���B��,B� (M���H�VVF}��p� �Xa�8��H��KZչ���J�� ��m�!�d�S!� �k�,��7�Z)�l(�7n\Du�?�al�b�b���,K�+��������y
�M�L�2{uzb��� ��t���r_�ɟޟ� W'8_�f�ӌ�Zd)}�qT���\+f��?���<x�~�(��[0-��_����e��T,q\շ����c�_���k�ݯ�h���e[�y�)E�n �e��!�x�������k����ق�[OZ�<)�ۓ�7�]>*X�w���c���h0u����l7{��*m��>�S/8WW*��)��X�y
T)��9�%�}o4�ΑR8���e[�]��x�Eh�FA�`�;I�	��ߞ����E�2�.z&��.�b��9?��6���⯨gzU�^9�L�$8������^+0q����:� �kbR>���� �r�M��Kʔ��}
��篢��O���*{�����M�7i�;�����g-�z=xB�ǯ��?��K�IX���]S���Wf���Pɤ�Ҍ �{X0�U� Zs����u:�(c��iF:�6햋r����iM��u�[o����pP`V�R��c���TwI�Zd,pҘ>�jODf߇_s�e�!ґ{�m�$�4��G��`����l��Ɗ2�;Cd	�"�В��M��F�'ea��m�c�'����{r��P��&	���<��'d_�tҊ���Y��=�;�n\��O5���.t�y�\XO��z�����\8��8z��������Q�&lP�O)`��*_+���}�h�$�`�MNt�k`��l��z�7�f ����l��[����p,2R6)�������{*����k��
W&/��p͙� �Cyp���x���E�ި�(3^�(@i��b_Z�,��)2��z�[<g�x��`I)s�!�"�4�(��T���'\��j��=�\�Ǒy��1�t|ai*�n��4�?g��/�9�9�l\�E�
f�����)�
!�/�C���͆���n@�U#�C�����4���eA�ttQ쇂��5C�(��3Y�o�K� ʤUO������Ϥ�"M�4�tPJ����
α�~�SQ�.(mb��5�tc�6�����B1s�P��ǩEu0�'؞� ��i�Q
!%�'��=^ Zc�_��}�d��[�D��2����b`3���%����	�bU��8w���E_��o��z���>:��(Q��|��k4���|�@�4c�Ћ:�=rb��E4%��mo4��Us�OC����Z���Դ�/�nϱ3����r�Ԃ��:�:�DV�I@ب��w��լ���	3��}cQmO����O��ӷ��I��t��i�Oώ�W���2��q���l�QaI����}�7��^�}, �N�jF�=�iha��╸ه�#_�nqNV�u+��/�:�оp�p�(�,�׌��FG��横斦1���݂�6Ŋ����0�d�Q����p�@�v9C�i�bॲ���#7�����j�X��C�}m9�W@,Rڕ@1��XY꺰�G\rSLA�ǉ��:�#2�4�	҃�q �I�^�|��G�"a3]���hIѯ�ۢw�����_��/������p��ϟ����.ݲB�e�S��n[�1j��xm/3z�o�2�o�;LKƤ��8":4�D��_/��1�)��nک��̵3�a͆CH�Z����\���9��S6� )\��y�z��~��
�����W�j��x
�{W�},c�CL���������xa��	s�����&h�cJ	�q� ��#8e�cZ����b��qT�dh�&R��o��:����*��_}^�"�_㐚I��m��e Z(p�T���}��HX���,�/�I�d�������0Nv:8Ju�S(��Qx���P�|��FB�L$y<bҕ&����������c��G��	�| �g����DUa�=7w��l�9KŞ�ᦠ�v�ʈ7P����{¬>�&w�J��3lۏa>��HW��|�]����2���(gy1��o�wR׈۲B|�G]�/���v*^v��X~{�d�E��?�HOE�n1�����Yg���~�(���߀KN5G�Ѥ���dT��:�	c{;L��ҕƜ���Ek�����4�B}~/�΂�
��#�,]Vz�?��c1$4vrS}^��h�$�&��4��'�M����d���T/�(z���4+�nT��� �(�c����p��!��<LǍ�:�6e
R��tuu|������'�ɼ5��O�$�Z�1^hh��}������Jr|���S�p��쁫��b�aT��I���l��Ft�jKC,űȠ�A��F�>|_�f!�b�4�# �'T�N����^`����`���P�E��o�,�#��W�̅�j�)'��q�ަuҿÐw�; �W�Ѡ�?�N�W�{�J}�Xw_�+=�v�^����8RcI
Zڣӿ�&䷁��M��$��يݮ�K��y���Y���e��CsY���!�K�c�����tc�Cq疿��6װVP
`����Ă���~8�?��|_m�C7�
���+�2�dL�e~���@H�I&�Sě��ɍ:�3�E�ci��O
<��q���Ğ�cOv	k���6������i����Z=��8 }���س����smx7�Us����l-�2�QzTd{緋!�J��j�\	� ��K �ȈS���h���(	�q`Q�C�]����aXd)�5^zU8�����R{�x���s��>uH�U�(�9J���{�����'Đpѿi|K:C��՜o��;Sמ�:Q�8Y�x����B1�E�OYN��� �'e����sI8�]�B�3�P	���wc������u�2V҂��i��s��D	��T�E��?0Xi.�v�M�B�A���]�of0�9)��}�M���盈�8��G�1ά�����bA��~+A!�p�6C��7��֔��|��� �v;���Q�R+�.���cר�H���?q��#к�.,��ĝX�B�L��)G�4�x�U��d�F��C�ψ�������w�E�� �t����h��������`��~o�^��W`�/��%�6�[�F.��Io��yt��
��$Si���RA�M�l/��y�$w�"ߵ|�zs�R��;CiGC����$L�#��Q�h ]��`g�G*TT��%o�[��&�����p�1񝒈t gcNP(�X���a�}� $�!a�aО��ȯ�y圱�%���8��x{B���ND1Vw!�Y�����Kl�V��MA�]B�	[N���L�b�u�n؉]�5��L����`�
K�}�+yz���I�S`���_4�=�����8M8+�U_��
U���>{�1�߰<Nc�uZH%��!�)��2��ְ%�2����qν�"�5�/����C?x��Ŏ������ӈ%Pu0��t/>�
���Ԗ���^ZtrըӾ)V93�D�d|���~�د�7�M=��:䒯�&u���������<P�k��*��9�n�&kZ�2q�ܬ���&��Tq��!�0� ˇ4e�o��ܦ�]�=�T���8 ���h�P��߷�)b�+�V\��*y9� ���K��.V-��|�ZYޢ�_t���+�ӗ[!�ʄ�Z���x�ח��㴰I���lV���9�x�.�)<ݝu��9�s��L3u�r%��j�%��#Z�ϙ*��G4v'��-dhepf6�=3�.�u��z?�ֻq���.��D��|X���:8����ӵ�ARS���'��`9�O�gj4��^����	�a�^��M8����7�
��W�E�5H���p�Ə*�����E���Ϣk�&���\��B��U�&����z(�	Tz��儜��M�Yjۙ0TY��M��Ğ�_��qL�+K!��d�b{�{v���vz>�.C���cEPV�sr�
��W�+�|���r�mD-ÈX��ȑ <ͧƴpn��6I��p�\m��:�i���48"ږ=���\Bm=$��N��c�܍�m�Ql�[f�A�!D�Q�Kq[^8���2�	>���9�
�癒��%v?<��ٺ���CUS������?v����:�W���U�d�ٹ���`�䍈*xG2?:�p��e�B��w[�FK�(�e��b��W+~��i��Y���d�5c�r��d�.���/v��@hŷ��r�E��X�
a�X��1������Xv��m>�{�0V�ɧ'�rS���]<�w.�V}v�$ �f�˴� U۶��l&J���/C8a�AHyf)0��t=ѷQ⑩��4h��9������8w �����r���p�h�
��w�O�l�|�vR�賕�{Jq7%+I���c0�.�)p����[��kd{6��7���VQF![�cD���%_a����m�"0�Z����B='��2z�R���/fs� �(�ˮ�LP���N@�6�Kf9'�/����ͲH �<��ס�~lX��f��%�H�}3�y�n�j=��T�I+l�A*�8Bk�߃�&21l'���6����pm>}M�)s
Yq�q&�}�����'J4��B�r}1� -���z�&%���䏀n�"��X��0��zKC̋�����40p�}��8xZ�/1�~a)���x�����ʹ�r�{\���2�w��]e�ɍ�"<��/6>�P.�L>��n鰖���^E֘0c��Aj���5��Gs����xZpԪΞ开Z����7�%�f���-@NMBߓո ͅSt XaV�2���<�Q!�ho�k���g�3�P���H(\+�R�gD!�*R�o���N5��)^T�6��l?�(0`�,t�/�~R:�~���gcj��A����;�T��Ҋ�4_F��Ձ�Gĝ�\."z2�䱘�����	s"
0z��Y��c�������P���Cr�����A�9N�����|�!�|���s���T����C� eZ���W;RX��2�QvN�ѡ�V��UeZ��L<�E�vA�����m�?<9��}C�[����y��S��fC��,�%��Q��v�,W?�^������������}�Hy1�~-Y�	��c]
Z4��&~��f��%�\NC��!�Jv�5�
��KQ)E���-�[�+�Vc�R�K!@I�n7E�$,�s7yՍl��&���?&pF�;7�E��[Z)��#�o��+6�)��\��()�s.:�`f6�j�ag�# �^���⸇T���tTZ�o�E�;Ɯ����x���A��|A�by���U�Vz
_D;<���r��N%�M�Z�C���K�5�_�L�hsZ��ȍ��谭��`�k��>��)Иʭ�g^?G��b?��5�w|�$3�Dz<��t��kO��G��U&��z����z�_ʸV>�h�@�#�6���`��|P$��G���_d�۩Nl�3������ , ����i2:iȭ(G:r�_h�2g�r��^��農��D�	���,��ka���e�K
��%��3X�g�"4~OQ��&鈔�R��2�W�c}R�H��5mS�ۖ�/C���t��d��}�V���<�,S���羏��K��!؂�Y2M3��u�t��XBq�8��)���Zx�e�v[BM6�ߨ�1�^�g�c���j3��K7�Z�2x�R�3ɏ��U��7��u�
�q?*i���5����vU�9��A,M]!�s<�=
H9���F^[nhK����w�g��*���n{�ȋBbz�:�q���]J�W�B��]Ř4�����\cұ�U߬�w�T�'}�S��av�Sʃ�ٵZn
M17�mA2����D �f��V��p�0�{p�&Y�G�
�>��=���mP�c��I�͆1P�L��zS�e�S������g�vsA2�V�����8�)�dٟnI��$ÊII��C(��	�&�z�1ty��[	V�hn�� B������[S�L�vL��^�(RD�KS@�	��b�'3��3�0�Y��3���;`��L�4X<*��lӐΘ�.sG�jѠz�����C?����$z��}^L3�qH��Fc�{�Fg�}��Χb�L�������5�����FLӅ�~��	�e͸_Q����O�ؿmvZ?�>�ڴV5���7�`{���H�!�D�ۄJ$��R��K9
�(�t�&�vk�������N��p���#^ʟ%<�������U`Ǹ�l��7�d��GN�Q)P@v����S �Lr�62x�T4�V�B̢��ͧ�D�g������PJ)"������.��ǎ�1������ׂ��0r�_��ףi�n��2��x�6}iui��wM1����ōќ� g!�īh2�!���>�b΋o%n�>��n^'��@Xe*�X����p���}I&���v/Th�R��V���`�kx&y#�Ǉ�����7&�'�nǱ.yZ��7jp�I�|�G����I�ؠP�eNx�2�(\7��pk`������-��"���V�� H����]�e��Z�ς��C�!cd�M��H[�^&<��B�F\�T-�ϲ*5�w0ג#��8��M���R�7��6v��j�1'$��._�JQMT֫�����`��k�����cn�5�SH[�S_�����LYib7�KuX����+�C��+�(P�5e�o���� 
��>�R��u�K]J�%ꗃ��H��˵��s�� �f�9�j�/��p�G��K���>/A@��*�THP2�PA�4��zv�q��w��J�	��T!�=#7:`�������Ω�R�F��Ё���&�Ա�`4�n���J�^s�%ߘ^e�$�K6Ṝ6#h�)��ձ߯���j�zx��X=�X��\�h~Cָ�z�NT�/('���%+J�B!��L��H�p���H;R�H&[�����H����޿���	M�l���P������ u�����ǁu)���'C��6���_�J����bdq&w��}�c:0��xv1����,]�� �����L$���t �͕�K�"$.L����Vm��5����;sb�ω�u<�t��ރ�޽i�t����s2rl������^��J��v[���) �qD!�ի*�ui{!z�`�Ջj_�;�l��P�#�Udo-b�8���a�m�wPn�-���\����#�c<�i�k�/_Ô�I�F��Y�*��}K)���Z�ϓ�q ��h����P;�4�G�B˾��3}�B>�@R���]}��Y��N ?���;]+#��}�W$�oJi���l��[�U�I`�����+�Tkqcǅ֙�C$F��"Cp��HɴtK7��i<B{��Ƿ3i�=��)���pyv�I�@I�?ރ�eNK�f���y�U��z���9ꑗb��ݘw�^a���z\����Ӓnh�֛@��Yu�mɱ�� ~ۦ��C� ���o����F#�����5&�*Dq�Ŧ%���}́��>s��I�����t3y,���I�݂��X(��(�ԣ��S�u(Ͻ�d��Zi��%���V=~|bys���@a��[��T@沮<��C�T�L�m�#n�9�R�+�}�I7;��L���&�D"?����R�-)Ix))�Rp2"���6�m���N�%�Ҍб{�:��0\�Y�[;1�;x��߭�'�R��V+��&~:����o:�G.����`׿;�G�x�9t�ړj����,�b��8�| [���q%� l�dhN$oI?�����i�2>װ�M;'���[���,���� �$�κ<9M�c�o<�8O�B�,p&�]�|�pᘂ��X.1!�����rj�7� �/��C������ohA�qHW%%����K�s�^=������HRm�R/'�>s�����zl�I��jW�����H-|,#����b�t��T���6.n���*-����
0�����s����л����t�2�E�-!	LI��8y�y ��\۽g�t)d�zĊ�ˎ��ʝX���6惤�hq"W��(��g�������P�����է����G�wK1�F*=�\����#�%P�7NԵ�T'��q�NB��M������%���<0��拠�P��W�^�>#���*�s�A�A5�&�|��A~�ͣ�2��"�<�@�^�i-{xH���Ҧ*�F\j�Ԕ]>@�q�d�Y�l�;��B�"9B�۱���x�VE��$���I��/g��cT��V�"$]G~�r��.���g�B
�������	�V&?ы�#^1܅��([l�5�b,HbID ������̴�����A&��z��ep�;�4�x>sk�m���jkT��m�ZL�& HM0<�P�EO[q�@U����8to�:�������C:��R��`�"���w(~�p%��=���!�Dg9�6��#Fh�������nUP���j��%����Oj��s��%l,�>ebֳ���Jć���vaJc��/��f�B��?���n��tz�"�g�]�l�"(��H��;��=��>�+N<0�޹D.��<]@�H�|v���ۓT���4��  ���+��*�:��'*[�����%��:��<-�;{ߏ!���H	�N���*w�Æ>Q�M�D���	+��|O
�=�D�]��.zp�f�W��J��VOh���I����z�_�������0��>q��'��I�B �{���y�~G�-�&"�m��d�c�LjGQc���������,�pı\������"�zG���Xeo����'��t:���דJ��7�ѭ��x|���c�sx��(�a{j?8C�1��|�Q����o�ΐ��>�v�zo�FMʽ6�]�'簳��v(u�� 3��)Qs�ؽpؼ#��r;9b�?%	��h����+XH�f��!�6T1^�U���f���A�-�2�]�k�*F� l'�L;:�e���A��a��6x�C;�R{�i��6��Av� 7)��6�ֹe�ީ ���@��G��?8�o	'�JQ%����*���6�	Ё�c�K��Dw�2!M��̓覕k���!�ȌE���ާ�u�qV�>|���2����rw� �!	5\QS���Z˸/������U��Z��߼�PJ!Uu��ީ�/&}��6��瞜�d\P;��9����3��xӑ{�kpQB�`hG�� yetG��8Qy<�˸'}���,mý�H����儃�C��W��V$�)��t����V���7������<U�ĝ zd��3�lo�Z���(U�F�I����@��^ϰ��J�y��E���`���4��<CpEz��i`���l	��+��ފ5 gǓ�v?M��k�,DETP�ǋ��ؒ�,d�8-5�A�g��+$���?�������dx�ߙH������6��T	���8�@^�#JK!Q����������2�OɄ'��@�4�����>d� f���..�5{H��5�_���ü���J �BiALz���^�^��|L@����}A)r�@��E��U���f�7t��5d�	�����xsǁ��-�{��i�;*+����|���.�Vt���u�!�֤|� Vb(�LLq˯���TV�HQ,
��kP7d��Ϛ�G�Hڏ]�f�Ĉ��h�l�~cA�9���T	6<������pi"��&�(ywF��)� g�HobQ(��Ʌa�ԅ�`��'��I�T�N�\�>x�'z���Z���Gm%@+v1��N�-�nѫk2��b����>������ [E=cg��������Ա~fH�v'�������
�-4U��*�V�tJ#ɉƛ��0(4�2���)����"HFQ']�HO����9����j'�Xq�3�:$hZ�f�-�Dh!^
f�=D�Or��˔
]p�G��R!�D���M���t��D*�Ye�p�d��E(¿�	���Ei�f�iJ�_!����~�)/���a�#����?�P�]K����u��y��w?�>���Wi ��.��`�k��TLA�,���S-lm��*͑����Ys��n�	�S��B��99�e�G'�!�
�imA�$��g#����D�.E"��Z��ZL|�� �����M��u��Ъ�oi���v���gr��^���f�D�h�=���x�-�i_{�1@qQ��o��"<�#�p�M{�芎w�_ J?��<]�������ғ�G��]s�|:\V.��-�j�H%�=���>L���w��9v�9*��m�݁$����������m*����f)H@��h����D�ĳ����Y�1����f���F��.@���U�By�~l��7�n��	�mHV1~'?<�/Y�,7����0ӎ�{L�3R�ap�׮���*�O�u]�,�К�K�����P ��C.��aSHG�����/�ʃ���Cg=4~��{D�6���18I�Շ���
ƌ����߆�o�]Y�.�L�L::��)�4�4<8��F}'ǫ��ܜ^ں\��nZf���5�0+�})P�^�̙�����:f�uɒ����{�S���K��HX�d���5q)���0�H����ԒƯ��n̱3%ל	��Qi<7	kSB{�v̝݆�NQ�s�3�D#Te���p�I�	��(S9�gb;�@�"[�� ��m�{����1��0*��V�&�o��H!��g@g��h)o���h��x�I|H���&��%`�����ذ>����:HDD�d
�!'n���E�)��Ԉ��"6�B�tyvai������#k��b	���� Ty`w�dҐ�������՘3�X�F��<�,�Y4
��|�9�l|�EE�Q�ֺY���ra�o�3���)ӄTev�-^7NO�)v�i�W��R�+y�W�T�0�5j�xs�\��k�h��E�����I\�P����`����"Cy7g� �v�:�5A�V�&�\��j��{��������L�����J�sp�Ցml��O�bn�y l����o�hE�?M&��d(�`N4i6>U��f72]�(w،�d]�ٔ��%ʨ?KP���ą��FY<���ё�ULB�ucik 4�~�+\`���y�/ӹ�+{��TZ�V$	U�>��ƅ!��}}A������H��V��p�7�U����=N���[��sW:p*'�[N�W�2��JBk��1���SN�f˅v$k�����K rp�޲^�����<	�'��H�:7�s�8OY�;�8��nQs�E�R򧥼Q4��[$�:���HU���wl���4�g(�/ܔ���t��s��V��{��I|m �Ñ����L��{՜�RG/T��ɶ�-}��~�&Ɋ�3K岔ɸ��3~@���6�_�	��n�v�4M����*FdSPQׯꗈ:_��|�]<3�n�@��q�xq+#G�MZ� ���m�	B, ��c�Џ�2�k��{��BIF�2�F����6���q��>�3�}���
Ǡ�h������O]D_�����)��`R�`v셱�x�l~�'��dmB}{cvP��o	6ǭ(�d�gχW�ݖ9����Z�RirH�>UsB6��Þ`��.:�Â�	c�\MJ��3���\������M��e��H�86J�����;��M4�)�, J��55�pv��i�Gt5��T�?��k�T�-���Fc�?�ܫ��A�5dlSp��9xy9� �ʂU���(���z�د�J��5�{��!�.u.z]�p�Κݣ�;��r�{[�<�l;P��'��\�Sn��<�u+H�/��zt+jo~���1!��#6�$�gjb�Q
��O��-PȲ���J�8K��ah����hA�(;�g��.�O��9=����n�}��*ͦ �Vz_Ѩ/�m�M�a0������q���l'�$vbuQ��VR~��P���<�^�|xE(��lĖt0�����8��{�S��׀�&Գ-nG�Ǳ	FB���cD�w���\�yY�����2
���T�Z��,�̓p�X(�k]�����lfz
�VxY��	-^10R�0t*�'߸F��D���쇪�mbw�6�=l��0��9褲�:�ǫ1�uf)�_��u;��F��C�����Gs����:A3Q��ba�M8e?b�b���Ör�)Ϡ2���P��1c)�,R���Ѷl��wY���C9�Xk%�Rc�������P�߾��}Y��\>�\[tm���$���f=����� r�LJ���@�x l���TY|b]�������f��y�L�ԉ�P� �9.�#N��)��=��P�����d��^{�*KC�2�UQH_]ڙ��gn�0��)v���o,�9{g1[?�� ��8���ҍ��}Q���Y�3�}��v��/�|I)�l�=O>%�Yd>�E������'|�٧�cj��q\1�p�E�� �]����̤���k���Xq��`�V����)�I'�ʀW��pc���;���ɏ=��-����>c�+O�=�6-(\K�aҐQ6Z�a��y��;�8>���S��6��0�$�B��!�.q�λ!�Hr��<%v��%��;�m	��gz���I�����{o�&��c�뢜��e-�u��-φ'�Al%��rsvTg�-���9�w��$�� ��*@g4�fV����XG�aZC���h�0m=ȧū>�o�e��-���M�T�.K]k�	��]x��'��2U��:��27����8��-���YAw� ����ӨJ,���X��O�0x�rE/�xQ���"�f��fdO^���t�x�8ӥ�ʠ��<��5ף�EM��ب�U]{.���Y���n5�hT�}O2 =����Òᡆ�����C.�EJ��g�P���X����3Oc7w4��a~{�ZB�q��`G_��5k*�L�qaA5�����{��eT��\���rb٥��wwg<�$B��L����%�zc��7E�fX�]nk��`N�V����<�ǉ���m�Xz�5"G�k0��&,�k�A�\!~)����}��3�[��b1S�-Å�,�vF]4�7���`�o��#~\�m��^���u-�CVF)1�tmI1��OQ�`;ƣM2K�|��/<|�a(�����A�����&\9_�� t��Ϧ2��iN<"S�I2Lx}<i@382c�%�S�%�|��,A��a�Jɀ^%>`��O5��L�:T��e��>�a��4���QyK/�����|B�I"��'��0~�c�=�>	���>;���6$�#��r����0^#W���1��g���E\����iL4��/����G_��#"�U�.'�)��N{,�m-�)|�mOFp�wa�iLwl޵LH� ʔ��P��Q�*Q�{)Tia�j"yᑉ*Ȑ����&�A0F��}��rb��&[Q���y���Y���Q��~p���t9����u�d<�)0�h",H��X1:����9���y�_8�����[�Wm���5��M����ћ���,��'i�6i	�e��o�ȝuA����PV�����4v�4�� ���;i%��'�O�WM�yy7ʝ+�2�9D[m��nlc�uA�ʮŔX�N}�8p���I���79�-���٘�`�ɽ�a]S_D2�_=�`1�M�S;�(+��1!��ӱPV[�V��@z�ss��l,厤�d��C-bz��HRݑo���ٝF��#�����E���8����p�A�W�^!2��C�ZY1�}��p�iݷ�Y�D�bO����ʢ��JVjy��x�J���yAꇬ�����G6֍�	�7�ޭ�k�5h�
%�l���T6a����xG1aU��s>I�'ŕ������+Vva]U��I�Y
�.25
�u�ù0?1-��!��]"��B
u�r���g� ㎍�G���v˕r�h�MF��!l;	�֧�9�?>�tuC"��w���x[�ը�����L���ߔ��V�/k�9�Co�1�q����.:l��y�-䗼\�q(��,��\sF/O)@�u���5x��=�B���/��W}x0p����Bp��L�T�h_��Lb�o���	�'��z|���^~��][n�M�����e�OPȿk'v	��;���a�P�85�Ч�:dZ�ͥ����ùn}������	�N�r/78S������v���V���L�x/=�vkE��0�U>�N\�L5�."T�ʹz �T��\[�����w�%�S��.ᰏ�l�b�h�H���Rǒ��j���te��m +6�2��r���$c{唲��w6-G��f�Us����+�B�7�J��>�x����K~2=�iaC\���>�`X�χ����po�WY0Z�""e�7l��$d@�8�6=�w�W���E�c[��U�L�w��X�����^��2�����C1����?w��WS�Wɥ�MX'wfܬd�����F�6��#��Z����7]~"D���֍����]Oe�
i��G&���ewx/�:�[��Rs�g�d��=�/̈́u�2e��m�X�K�a� *��1�_����i��	~t�d��X�ߡ�/���V�Т�����Z�,ʳYnh1�H�q$�N�B:��归,G)U���Gl�d�hw� &�E�7id���j���ϼ��!ݩ�8_�q*E�P��!<d҅������{��߁�>m�xL����?{|66�m;�������7��F��ճ����8��-�6N>	����{ƒxE�#y1?��#����|ȬdMjǨ]�����TͽML������=�*l�5`��~��}hz���0s�5���^d����d��g�/�Xޕ���L_�U�����Ɛ�����@��+���_���A�q\�dk�|�B�=��-A�~���-	��P��#�0�&��,{H��$�4
��p��`ʀ�V��K��?�Z��D�%�o��>8�՛M��e�Hp�����gMӨ '�.���'�iPe#!�Q��?�K�s�!�N�Ҳl��t힋���p�hbk��Se{�Q�8�k5Iʊ������M��(���@����8
U��\�G>����-���^+�U�bX�<>�N>��Nvn ��P]�������D-�-����=��z�g_|�hGHMM�n��BԒ�1w��#z�ׄ�W��i3,���G�3AK��~���2�şƴ_�H�n���[?YK���7EݟF�SA�	�.�*���m�����jX6��[��Bt0�����A�B9�(��-_p�]L_�g���6Xv"��� �ͦ��J��&�K�Mwr1f4��|�.N�倹���A�YA:~�ʿ_���d�	������g��u��7�/��s0a��r�71�G�[�#�_�Dɇ��ъ��;f\���[����n|����.1q�D�H�W���^0�^:0��r��~��Aߢ���`��Ģ��/kx8�u�D����Lx��̪��ƳA�� �_{��Y��,uC�m�L���G�c����5dNFb�0,��b��t&N~f,7v�&�w��{&y�W�o	�9+��VܔP�*���$DWX��Ρ��z�*���g.2�n\�mV�v�c�P���d�u2��1��K������=�X��=�P$��Q_�����Iě>P�4
�#�����P'�Ø߹�%�T80�����P�s��PKBm�$�kٶ��
��&7S�sS�틞c%5�B�8c�"w�cN���Q��E�&&j���W5�m�����_�B��dl��M$-qF�;zR ��+���'5�N�$�Մ�9�kF�F�v�D��J���Bʣ�\�7����A^���Dv	n��D%׬ن�Af��j�St�Q5�]��b�B⟨�;�Vi�`�Z��bC��j��cK$�<���'b�e�K>���s�ۖ��?ks[�k� 
�1%�@����� ��	|N^��}�4H�3�W"�^�ߙ<�W�(��|"if��vS��̤�7a�mxL��I�{_���A����*��	�k�jc��;!�m�uE�����O�@���&��,�
�훜��,��O��zE�
 1��ǂ��;T̫s�#���5��x	'��G/	�3��jF^�t�/����ݼL����ĢX�ô�ټ6��֧�SQ�j�pl�:��5�bu�,QЧ��Aۤ�0 �6�'=Q
��G�a&م%��J(����"���$���7��+�|$>�j�͉<ҧ<��k�ݘ4������@����͌��|�T_��v*�;r��\藟�Ww<Z��%B*�~��	�+�p}���9Fo���D*.C&��A���&T~�ׯ� �m_e\�1hCH mE�_��(�(�.���r �+�:`�IC�o�ߡ��@���"h��J�v��h��J2�50�Z�;C��r����6��E�.��Y<ٲ$�h�//N˱�����D���r�N_0�b���A#�����=-����u��|�M�A0m��/�D���y�0_1[�о���Z�5=��>��������U�N�^�D=�m��q	[����x*�J�Us�k~��%���$�;�v)�=E(���[��O#��g(�a�G����䗕��tvQz�h,Ȣv���*���;�@�1C���i��W��7԰�/�>����
����8Jx�ɮ��~
�.���(�F��1j��ˎC(9Y�*�������[�Ԡ��,/��KLl}����6.���on#��D�5Y4T�ǂ]�	�0���_�G�B���D��$���3�	��v��t�[��/��H&���2��^��
�ڄ�/AE3�C��z�[\2�3q��̯�kl}jp�e�*c�h(b��L=��H��p�����Gp<aFP,�e]�s������rHr.�1��Z��j�=�69�p�\��ţZ	��~��$	����&�X������y�&�� L=�	]^}�Ex�b#a��s��f�!T�&�vy	J
Ev�Ἰ�^��<%�q�+=��_79m����?��(?��f�q�Qu|���uN(1�a��L�ͳO�h��UX6�b��m(%��Wh�c��mF�P�AF����-���a�aEɌ�1��юԆdXJ�pW���}
� ����P��U�#���.9��v��j$��1��6��)R$�~H5��N�U�7G�C����Lؗ���K�1����UH�K�\׻��S�{1?^��P��/�����
m��ɉ���
�<��
�N5|\����M������-��X)5��h�h�Z��.��a�<D!uÕ��Au���>�i�k'�'
�Fmk��6M^�5��
�-�c/>��Y���W�Gg	B|�L4������ճ#���zPJ�b������Sz=�Č�0j����vV,�a���|�,� *u���N�B�Ƭ�<(#�>��2���֚b��!�߷�~Ǣ4��#?�k�T�)�i=(�ˋ(��!7�I��j,D��i�g�VU|f�8gZrt�o�3v;*L���y
���Ѣw��m��n�o��^~���`ξa��
4c�;��%
҇���4	��!���5`�3�h����ԗ��a.�|�qm�jj��h'�gӣ����Y6D�w�������K�]V��F&=��6��n��>�̂�|@\��'v����N����
�Uc�d>�T��r��[<��M���A��b�!
1g�"� ���TG��sВ�3���!��\F�ӓ�U�BTd|��S#�_�Ԛ��K�õwC?�:��VMc�8�eR}l�BM��#<ސ��D��*��@W�Ag�*���8b���<��g/"���Q��K�,L�Zv\U�W,y1m�������B�2����1��~��u�7��s�G)��`�萨�i�푆eq�?[�%���Ko���]{�2o�%L���r�	Y+�r�P.}�\���D�g���;�
�ݾ�I[��J��V�O��!��P�#��q�c�c�T2B�PT��Ӂ��*^�'Z�y;�&b�)���n�����ɳ��OK�,>]�������B��tќ�4WSZˬ_��S��ӾK*���@�U��1,�&G�U'�E`�����������$��y��:�k0��2���[�g�?�Aӽ��
�����{
Xx�]�!;7����j��[10�m�Ƙ�e1��J�����i-t�c��ζ�3���N-#'8�gk�]�aS �0Xon(q\����`�m�� ���=���n8���Œ�gdEد"�/�rD9��\+��.�x�F����!�Հ����#����(m��{g���9�-W6��mE�~<�Tvlb0:�uz��$}~��n|nJ�h�.f�yj�A�d�y�~g��sf��A���z��`#M�Κ,ă��zG������C��S�=!E��LO�qZ_����B�1�"�mk/�gmk��T��8�`�%/bw�<y[/`ڭ�Y켰8��|n��{v�@�a:�x����u����I#rp�#X������^?����<І��	p�¾:�Co��[}�ے$H6�o�}�H�F�0�qr�P����k�+��p��|e(D��DZ�l	-;dl����j�ip�@&�v8RK?�����?��>
���<��
a4T�)ڜ�ױS��[\� ��� y���\��nxy�F�zC1+�Ǻ� ��D+�^�r�#@��,:q�!>w�
(	F[��@�F��zk����kc��?�o̥N{�2�8�{�#�H0�^ո�|%h�����yiJmV�ԟL�5�V���_7uf/���V5؟m��>�'�܂ؖĀY��o4����H����rH��̆}�j�1f����F\��T��j��<`v��-+Y�7��k+��7L���Ϫ��������.��ٹ�!������@pJ˾�
L7/�R��G�QǍd��눙$������$��,'s�-���?N�&���V^����^���A\F���	���m��P�7k�YRHeZ�Y�i� �3�a�hD��˻+ǽ�n:>�d��,j���ޥ��US�BS�
k�cY��U�D3GWH��b;4�y��h�!f�Ye���Tv��p���fEo�������n�ޮ)���LASp����b,�v��ng��Q��������pn�����d(��37�Fl
�,����JHr��Co�c'XMD����f�hZ>V4�)��H	�hG&��:�#��.W-濆�<��d�3ɷP3��.Uzfw��Aݷ;�lv�H�IVUO�
1�n�Dc��5t�	q����v~�����T�r�!`�O�4<~h� �+`٦Ɔ� �Y�:Pgl
�'��~�XG��$�`���L{����pZ��hR	�<qr��MQ-�5sEc��Ȗ\f�"|�2��>ހ������N=(,^6/M�aH��e~lx.U�8[� @y�gBЬ`<�F�_�֔� o�LK��Z��A`����EĻ̚��a�X��4�S>��I~ɴ��y��H��$�h�@* M]v:�Gi�' ;��uέq�!lځh� �Z��bM�e�$M�2EdwyP:� <)��_���p�;��
��ݷ�E�aI�ٱd
��-�Îco�D6��l+��gcRc�r�<��P��\~��:%8^v�[a6/���Z��ɸ>�=rn�e�|_Mj��+��Ck�|T-�f�`�P�cgv��v����X��2�:Q-"1�Tk�A)�� �,���ԮWJA�KRoU�&�����vzv�9�x�YW�g�������<`����)�T[^�n�1���8F�w5��u�͏~�������{��Ѫ+'ע[?>'P��r��� �R1�/�C��X�mН"����ٛS���<D�����FҔ�C�m?^� }�5=��4�?�����C���UT�y��I���d�yq�UH�J�~�;��[%�ZD�^�'Xڣݽ�d;lmol��f��#�S��31(�x��:ǹn�_�>F4�~M�&~n�&��w,�/��U.᫐`&4(㷐{c)�.e˝/��<mb�C����c�����`m�$f���P9�����#]Q~NpG[驦�!� M��5��.ŕ-�V�F��b����L	��vi�<R-�w$f�YO|�#�#�a�*����p�U�pKޚ��m�İ���boh��b��1޸��$ 1��V>��DB�;��x�%%�5ҽ#���N�����TņToo\ތ{'�L���L�+
��^�7>&�,+�Dx�� �m'�A���	������G�Ϛ
W�b�;��{sܕt�T~��!���#���JXo���yf�w=�*������4��=L/���<�y���w��0@���sw((�(FT��5��K.Ͷǆ �܅qi+�SK�4K��0 SB79Z�514Ǫڟ0�[RYW<ԁPD��K�R8�
���d�`:�����w��(c!�p���N��l���D�����YY|�"*�+�Ә�Q���r�YH��&�釾:��ƪV�r��yQn�k7`"�>�i�d�]0q͂Ems�XXY��D������	������ 6r]��0Fܕa	9����h�o<�1F�J!�1�����U�7�������V����# �Q%��+a��3�ί(���>	K�5P=3ӶC��N|`F�d�Y��5�`<F��Z,�G�KUUw)��KlG(��*__���\���|xEDҷ��$�fp̤�Q0���d w��I�r^��_(��Ӈ FsI]%���|]�h��/߶�Oevw�����뙛�b���+t��2??�m��^�:�U	͗`���Ɨ튌���-gE������܊tc�E3q�|@�ߓ��_6K��3�
�jT�d�P	 z�LY���O5���
�z��fo�t��yM���A�`�q:��A��:�o��fjn3n�4a���'�����C��v5�:n�;�y3�s�\�J[���D�O�SA'�5$�G�Q�qm��N��PhZh7��[I�w�K��h		�0�%��D�F�-��-��=����p�����`[�v���.���ti�bO�M�T�����m���@�d8����~��"���:��GͲT��|���R7=?`]9�(�6/e���'@�'wԍQ�U�Rk���D����"�	a���"�����L�Ia����;`�%-�Е91d�ZH��q1,���������AL�\k'��<��E����9����E�wq�!̽�#�ŁE��Ʒ�J<��N���g��K��������	\�0���uբ�_~ܾ�q:���'?s`��ex��.��ƑR�Ml�y֕c��U,H>׌X���P�{�K��t��?$����L�>7߶H��	7	�����_�n�"���g=��N��\�`�ΐC<�˒X�,�}�FԫYL��Hmvp�= �F�6nP���ه��Z�~N��؇�--%�������[�W�f�gM)�""�,�+�ݜ:U}���O �)U�>�W7q�e��Q�j�Ba5E~�`�?!S���q¥^q�9�5�}����!�(��i�Qj=�S�x�N;���0⠗�Y<<��Ж������!��]̸�h��tx(vE
Q ���%[��� �� �F{���	��6�ʹA�f�c\KzL����=�Ŋ�5���������ln�r֌��[Q{a�,.mD���Bu�p�W��>�{%��l���U+C=$�X&��}"��8�k�.�I?���L�f��B�TФg�U�<��/I�>ւl�^����O��,�:�f�J�ceg��ڟ%��ji7舿��O��d||	���m !����]~�({�+go�9��-�ƫ�Dn�%�yɄi���T�Tr]�rN÷PL��
:?>�}Q��{J�S%����f����1w^��`-X%U�!՜�t_]1+}4����iHRp����ד}�D �Ź��[8GG���P]��7��z���Y1&�jt:�?.�хq�u��V� |Z����cP�o��t�F��� �]�nM�=���Ӹ&���Ϧ��d�"f�C$�POVb#o$06<�.04���%u҉:�ߍ�w3������xﱙT��?���W%��=�GA�����U��ë(qC�D	up���T�i�+TL�?1v��R��72����������Rb���q�Md3ɒ६��wK��*���<N�D@Dq��	gǎ�i?a�>ށ磽���h��^K�b�ކ5��}j3̧_@��5���V�\��%['0p��ƥ���쿙}��X�N���<M_�X�`�8u�Q�l�U��1����N�S�-x�����*�զV���Ag��h�h��W�Z��V��Z�CE�����>��X�Z�%��ѕu�`��	�*ol�hi��L���Jk���y�a!'�bk���p�4�a%��Y�r�f&�+=!�QA������Y��\H��V��d����8O�!p�����ɬ��WC�E���i�2�#��Z��F�&�G6�B2�!���DX���ےf�oP:Y3���/ԙ|��O1����iI�wʟ��{W1�Oj���P%O� �ќ��{��o�,�|^�Ik� �;<���z+$��%�f�c'�R]���m�9��J���C��9����NL�-��)4UL/G�D����+��a��#B�!{��V�w,A�H��F�Xc��~������I����h{���f�]�[�2���J���#�Dݳz��c.B]#����țlp��Kw�`��� q�)������zl��G�� bzT��`
p��fy��% $�s��H<��}Q@���LMQW�]]����`+�V�b��Km���vҺ����sl�<����!���� �����`�V�?0:S3�d�G���;=`���7��/r�v���v}�:���yj����H��L��j�ی���0��$Q�)�����pOԅ"e*O��M���Ϩû�J��������Lf{.��~��4�&����8`.�\Q�|��xW��	a��}$"�?O�u���/4b�I�_)���}�s�g)�w"ĩO�L0��l<�h,K��ּ-�g|VI�����ZV[x3=��oϰ⟇#.E��7�Z�q&��l���}���P 7�&��X�f8���]�ꧺ��Z�k7Y�R.��ETf؃��A�ٝ��|(�z=K�/"��[y�pG���=?瑸�L4��H3����镭	C����Vy�']��l~#�Hc�I@��l�����MI��	_L,����s����z�@����~�<V-9�aK�V��	,ok ֦�[���^~h�麟i�m$ߓ�뉃B���/�����l��P[6o�P�r�7�p/��o?�(�?�\�Zj���k��������
̒�i�Xr �y V�-AČY�2O�Q�� �<���\"L�ȣI��z�PJ0M�J=��kfc6)��P�P�Jك�8�ȻO85Av�#�(�ْ���P�����;/�Od�0�9 e�B0���K��Ok_��76�4���H>�3&�<�۹߻*.Z!� f��lNZ���ѭ@��RQR?)7ò�nx��E,��?o�~�g@�f{�Uṗ劵\	�8r�:��.�q��q��������+@6�3��I�[Ҳ��3��#+g�K�=��
�0r{�c~.��cc����a��]ĆmZ}4l�j��9 4���l{4Z��
�M�)ћJE��?����E�^�%��y�����~�urm
����,4�
�7ʕ�"��v/1����w6�jڪ���M�����啒�<-��mn�ш��J�p����X,�-��eV�`MZ��X�[�~�c�Q��},��~u�O���K'�d�	o��;��G~��1�7��;�����(]�N�$�p]}��u��'m���?�r��2î�o����A�J�#P��i��'Wi5j;���P�m#"2'I��U��di@'H=�ݽF�)���܈�;xq�� ��v�^
����sHWi���z���I�ȝ�	r���^M��{?3�ݝ��xN��o`��Q�ǀ��l����Ml��L�HJFvE;�6��09� ���G�g�ߣ�"��Ż�Їş�����"������
�Xs뒌|�p��+O1�G��Q!��\�r�?���!Īh�AkOl�W���A<������@�J�B�2|���	(_z`�63 �+X�ʧܩaɭ�G�s���YӖ�p�)Ѳh_d:~����g6Ei��r~0�"*��8u$&������KJ�wL�V⫅��+�E4����e�r
L�R�w� Y]� ���|�!"q��0�
�s�E��%O %iɬn���Oda]��W�n�S�����S���8�-2����u:�.���o��{��2�p�u�|B�'
�$tU���awP�̀WL��Qr��<i�ւhj�' ���y��&��Ruҵ��Z�l`C�=S`��d����9�ю�I��;[yQ�0�΁T��NQr��ç	6�7����O"�8���\���'wh��M؋6 ��꺪���H�˹+K�o��!xe�:��C�I�'o�����;/I2�nQ���������)��@�9�����٘�v�u�u}c��o������E��p��!�]�c�r!�񟼷}Vi$�;r�M*a#ܤ��+���-}v>n�0��`n.�ޘ'ݪiQ�`ޟ�h�%8"�@It��fESg�~@t�"��n���y�eQ/9,0��?�F�v��UJ@��¬�A���q6�X�#@�����5�a
qu�I�<�?� �ۗ��/1$���d����.�I6��5 ��n�s�5�34@<4���(Dr.��xa�nn������Բ�M$51�6m�h(��Yq��yP���j�ܼ>�-�R_��3��V��OEIp`
�I&&hO���{�IћL�g�������-���	GI�J(+y
b����+�<Y��ǿ��6�I"�N�-}cA�6	�C{���aXrf�m�w�ivc@�o���'4K}"׊�:b ��}��6�~��R��d˿Y��'��t�2vY��6�s�
��S�v= ����&�������r>��#�W�a7��Z�e�O�5i����Kȃ����T&�õ��B:N�ᘈj���sЁ�;��QÂ����\�-D��y��\W�: L4C��iQ�����Gq1-�VTPBs<3�[������7I�t�o �ݯ�r�����'O�%�[�?�G���?}���	����{(*�"tfB(���C��h���F�$%�)�#�	���	o�G?
��q>�p��x|�Oˮ@�k{�A$zf�_���g��F�m�	������8�M��1�Ɩ�b�������cȂ�����\J�^�f�C^�{�~���4��2O�邘i䚖���<���| o�P��+>&/�7��Φ�ࢴ�f d�����sa��S�Ra ]�".�)���̳x?��
Z)�m~�1��i�z�U��A�cO'c�ث�Ȧ0i-��j��B� �c ́�廠��e�+܏v{����Sb^1$���:��������6�^�܁(�3'�I����֫a����ۂ���u�y�ݺv�>��@	:M����S��\ch}�����΀��<�+\v���{<D��v�<jh<#c�����ćp�n�8e�|��3���mz^����L���Xd��Ө)��O>?Y>|`u�Կiq���:�bi/(��ޠ�=:�_UaxA��l�_�k��جt��w�&�Eg�������'H:���E���� `;} 67��f�ϡ��g��C�L\_�,�ʌ�|B��P~h�- ���a��I/��5��ʢд�ԓ&�{j�-�n��l�\�k��61���:�LL%�X�� {\������ Xt�,ς���,x'z�1�S�	zG�dl#M�`�0lD��"���l���K���Đ�X���܇���V������9ֺ_׋�aAH�
�ǹ�*;+�gsٵ��u-�ǋ����;1��]v�l�-./�f�^/۔(٣�=@_�N��p����Y����Th<:^܁���zZY�%�/K[p$�*��^_���cE&���)/��a:c��8_������x2X�!_�)vv��Y��.����O�Cl<���/TUJ�<����������:�Z]m�Y�Ex\ɪb� �k�nP��QR�y&}�]Z��b4�z��s�}[����|�z��V'N�(��욣5���/D���%5�3:��X��8$�o��6�H�������&�,^ʸ+�~T�)���\�J�A�W��K�\:����b2_�.�D�W]�Kw	%>�DE*�}x�1F�y��`E�T����c9௿�g��+���l;3)ݧ6҃�YPAj�`A ���8��+<����KJ������%��(T�
>�A-���͸�~MQ�-����;�9W�l����m-���"��y� �o5��fG�M�RA����-�����騋"�&y��y�I������m�"%I�e4�S��ˉc��}w��J�י���=,� �1����Y���WՓ�d���m'*�����g?{��>�n*��!�M1Y8�۬;��M�i�1e�t,z��!oa�q��5��Y�lgݴ��lܴ��M[[�Y��X������^G��i��~���&�!5HQ7�1h+ލ��h��_v�������дh�*% ��`C���.��Y|��@����)�g|dPoYnu��3�W�o7�s�;�gB�+��/mȃ;&��ؼC�������E�'.�G-�	�&�C��cJ��~�d��p�{:_��?$`Y��Q��5R�]A��X%���I��F�5I�S�1��Ժ�3П���.a�xQ�����r��l�������h���(j���l]��g�֮dSI�)D2�	���s��|w�UB�Y�,K�W��j!{n<P�gwN�]hS��D<�D��h�n�En�>)��!���tzt�����hxGC젬DJ!����^3j"BZ� ZX��ЁB^���Y�8�+<2M�+(�V6�L=��q�@��a�E����M�(���6�$��� �~�EV���P����_�2��p�����pp��B����_iW�Xn�F�H21sX��p1��Ӭ������!�\	H]��V�n���|<�!ij<����F 1��&O�恣MT���#7�$o�����0M~	>�R=t��bk�s��J��zɦ��W���GG�Y���b],^)<�<RA7���܁�{U�X=��T��*��o�������JM�Y�h%�ҕ��9x��}��ԟ�m�uԾ���nNG�.Z^�hՇ�l: ����$oo��gk��K���&x�I>���ޡ������BY��������_2�2�'�y��T!��gi���~�����c�����~�}���syF�b~B����.��sue�~R"�U7y���|}_�\��~iQ�?��;�=�38-T<1�_]��ե>�,գ���#n�F�δ+Pwy�]���Bj�Tv��֚W�S �c����T����\�3[��H�}�8'���O݆�ˡ�xi���ǋ <�9���%!u=㳍K@D��(uX�X�$��$�˝-��?t@��\�*�*'��X�Y�	[D�Mi&�<-��0K�{�(��,��r��FCn{��X9'���,��0�z�*פ�ҽ=:f>0��F2�IIv������C״Ϋ��{�̚�i]��?�(j# ���!:�Ⓒ�D�U:c�	��;p����%�%!!~�~�q5[�(+{��
p!- A#'E��9��}�����]0鷓��~�_�R�)�h���9
�[ ���V�X���,���qq ���R ��}������e���X�47�׆Y�����n�.�(l,8l�����8����v�u�C��B�<���i� �|�c4NE�]�;��H~��>5���M/A24
S?p����kP��B�r����ԯ��gZ'��ybp�í{�;2�6rk�i0X���)ɸ��ʤ�Q�L�j��,O���Ȧckd8���P@��1��b�\��t0�w@�٥�d�H�KqV
���HfO$�c��ܯ�'�߱�9I�?p����3���n�3��dt���Y\� ���&��5�,;����#� LU ZS�w���d����#/&J���15�P��m��� v�c�G�F�!c��zoL)��=����I�C��Lӥ�����v��S���\@��w�����-.<�aIƜ<D�%r���g�0���|Ʒ
�P`Ԙ%Y�Z.�z�3�#���د�DɆ�7�h-{���A��o����0�*�q[���v$]&V�X?�������q���;����VrɦG��Hm�#N�S��J_��ݫQ����� ��R+B��L����� �4Gg������������͚�ܭ�P3E^��*�r��h�vt	�F_(����p��>�'O@{����;,"�������)fgX�Ƣ@��&��B�A=Q o���z��5�����Wy��u�^���~��]#ެ���
�ጺc�ދ��@0ns�id}z���ߩ�V����£mw/�sde���f�����}>��c�����@��X�h"Q.]e#d�����4�i��շ�\50�	"\A�P�2h�yڇ!�����S�\�f��Ӫj�<t���YG�,���CR��:H���WO0� �L}�l3Jx�=���5����5U�l��=Kod�D�W��+.��<�;�E�@EU�K���7�i�fâ�Th������S#B��/���i��DR>���?�=ձ�#q�a8^M���k"�S)Mg�{��h�
L����X�_]n��ݩ
�2�|�������	�|Ǖ��+��Z���n����a�3@1���~��[2
 �:Y�[5`�Ϸ*�X&nax�؍I
T~�>:�c� ��U�P&Ɣ��jbO�'�(hI�8�7%�'_�E��獝`��=]�MGh6�;�
�p�%�7����e�Zn�S���Xx9�#�ľ�F�W��W�
j�"�D��>��?�#E�)�M�xl��ŊlS9�����;ڒܪφ�a~"��v�S��et��;����*�|=I���s�%��#C=)^���(��t:}xNl"{���=o>,��&?�p��oJ}=�V��Fv�~��A�<?���#"����u=�	r�����GJk"�O0/#�*h.�'���PA
q\J"=�viz*n_Ӡ�d�3�f�o�r
�ʡ��+������)���p���+�l%��z����T�S.�՗,)�P�o�P�Iy@���Y���� r/~�[zx��Pgb�o��l��*P��1�e�(4YVׅ��<.k����\?���K����ߌf��)�4~�������r���rT������P:smtg!�LGQϫ�D���^�����b���O�N��<Ś����B��t��\٧i�k���v6������6 ����K��1��8�ol��	1�/�z��.��֙����(�k�?�|�&@E���t�!�5p��g�E�+Պ��"��F⦒<E4��'>�����ft��S�R^F�7�J�h}E��}�棜2n;"�zo
c����.Ԗ�I�$�m2�u��r�s�A�[��+bܫ�I���&DZs�}��G-o~J.�����}.Hz�HJW�>�+x��F��3��s�!�	�xg�/8��k���W�Lp�������-�6�Z��7�[	WY��{x;P/�;��$��}���p�a7N���Q�EQ�K|$D�*�����FA��)���5,d�bo��O�V*�ѣq�U�{�P]�oY�xß�����	��C� ��Б����I�Z��]���^��N]w\g�"�=��1ڴǖdhX�5�1`c��V���25����!\���4k�϶�u0!�%�ރ"��1gK�Zy��2���ޜ�sD0P�sH~�g�'m��]o���f͋ ��g��niD'���0��}��/�����W����P��lF�e�)R�*/J,T5Ԅ!q�y�;�	k�8�!����vY���&�.+`���3iɭ�ϣ#���l���@!LHSó�%�Ȗ�� ξ�Hڂ*x6n�>�4�#�����m�Cf7����jQ^@���5h�����^��M�����З��X����-u��������|��4d���쭤@�*^N�1���ff��>Ѯ���hِ���<��`��r����_Yo�	�������y��Y��mR25��2��W!�URZ�.��6I��P#�a�`%ӵ���2L@M�~�IB����`u��r���3��ܠ��V{Aʏj��o�17A�ߞ���L�f�>��↳�~�	OC�A̱�[N:PcWN�Ew��Ѡi��
֬b����G�Q����E�����6���\����Tԧ\caHz~��~��G�I�zdd
����u�
���%׾���h�+sΔTOXE����{
��"�g@I���Wb$q�.d.ӝ�ȿN{�$T�y�]��?iTQ�y��A�V@.�/,Nd&���jƭR�2e�Ң��U�@�X�;�xa���8��leoO�D��6����C۵�I�򰊨K�=�����?}z���,�9z$��s2�!�a[0ދ�X0:V	M����wǽI2<Fj9 ������ WmK$HguBri5wM
��TR��bӣ��ۭE�ON�"?�=C���:�f�ʟ�3�0�M�����+��]qY����cj��#%|I��T��u��X�8y*�*BK��I\��ܝ�_p��h�yU����9���`?z_Ät�L�2��D����e�#��4bźglb�v����� _B�2չ��	tt���pF��}B��}�2aa�ڈiV�^��&��.:�
$�1(���s�3�)M/=|�}�Q�7U�d��_�v�QD0~@��k���K�|9�_�F�&��:��ANH�a�ŋU�q/��g���F$|+f7�I�#�H!�9E�=�����#[����[��E��Y�UD�̹2���ݎ��R�0$"/�rl����3�x�%�-AR�Ɖ�_)-���.�j+$�Xs�4Q�0XV�[�3i�#Y�\�qT�FuL�{����aN��d�u>u��x�r.��l8�Ҏcir��X39��M�`Q���-�7�2��#�A��#z@��8}� �u�|O{(C���ҋf�)3�QD�ᣳ�2WO]0[�}�f_>9Mġ�4~(�Y#g�<DޒŅy�3�k󶶮t�RT+.RD��0	'�r^rw�JP�a{�&v�����o.�!!���,5z������H�V��x�X�\���Yl�.�-~��l�9 ��q��r5����T�գ�׷F,��״��:�:�e�<&;EL�|���|%Z}&?�wn��[����0E��gX|�X.���Vb1�㾌c� �����j�h���AO�b�n0i 
|a�jW>Aä��Z������ȗ����B���18i��2g�fa�^ED^���Ɏ�]������	Z�#���ZA���uU�|3[h�������%�-/����R(�����L�)	q-i��A4�̯�1��j�����w^�
����,D�Yh�g�O�s��x�1�i�V�7�w)��$��ie`�~���%�R}l�Po�qH���lL�ހ��w��Q�ca�K� ���?��	�J��A�]�_��kw�uA+v���G�:8�����OviRv�e���f �릉��k�k޺
�㙾1Q*�"aƹ�Ӏ'7f�ٕ�t PCFU�����ka�x9���[MT�R�.w��N+-�J��O�>�B�l�o*Y0ጭ��B�]zE��I�M|L����֟�;o������o�M�g���U	zR`� �/�����Դ�l-�)�����l���5��)���wҋ>c��<��q^�@z�V~~���7a��7�yR������]��6{WЃk����ts(��l�j~�Ǌ�-m;&��"���P� ���:o�Y��&�����6����)_ٌ2�C�ǉo?���l��_��]O��fxSJ/>X�v-s�g����J�+M�Z����}^���J���͚ڝ
e���"��QO����W���p�[����!nf�R5-N�Z��UY�^7�r��P4�塃����LD/07���׻�Hh&y���"�rLE�߮���e���nB��9/ܩ�+�Ejh�Z�ڲ�����-�yh�C�X� I�i�eG~77H���u��՜���2�G�� 	��!6Y#Mz��)[[� [�����Vʵ�}�sk���u:!�[.7��B�:���b  uZ��jwH0���P�1���kGh�V�)n	���| �>���͎��ߊ�f^G�y7�>cˁ������PD��!��h�uv,�*�տџ�>����/]�S{���$�@������m��pF�Z�N���b�뺉�r��~���ޠW$դ�s,
&��������G�"��{w��r�s2���-/�Pն˘� �gC��v�V���Mد4G]D�v��I䷂�����*n�)�K,�S6^�"d2�N�&Y���ց���V��0o�~�!�U+'��yR��`���ԕ����R{��f2r8+�{�<��QNT/�+����+�I�=r��`ɦ)x�9�N���7<���_3P'GC�,��Z�a�C(�`�~,݄�v���������$�#�P+rtgO�(#߽������Fnc%��-�|M�T���G�t���`�"W�KgK��F]>�&$�s��t�F~�w{: :v�.ny�0
.�uLJR靼��D:te� �B�8lh�$�c4�CLj�p3y���r@��r�P�x��:�?�D�*�Q�i(��EV _�&7�$'}/}6���1�����1}��j�b<#y<�F�I��l�v��b��h΀��w[q����A�?�f�6����R��Q= �?=@Ŭpǡ�.�d���C;^���J��z�‬��\VO�hد.�AЕ�ӟ�;a�}�W��'��t�<�L
E`)LGJ�}%$�d���tZP�gT$d��{�S /0P�
n7�MʠVd%�K[� ��~�w�	@�񴫁�R��q�߲0��4�.uI?2�.�d�r �.��9 eS����9?�٧���wөo����Ӊg��@����ߡ�����9��}��!�9�jƛk�J�g� t�K���_H	�4�1�lDF�J��vP��ė�:�f1y��"�੾ƪ�tJ��:ɢ��_�L����Py�9˹I���CP!,����C�[l	u��M�k|�	Z�.sZ,�SZ�~�ˏw%����$2�gP�r5nC+��
W��&{���m�<,|[�k4��u����H�w
�u@ѓ1p��[�e�;*���[w��s�Xߦ�Q�uȪ;���`�����x0�N\��w��˚��Qo�P\�S����=�m��5�A�Ҩ�s��H'�����r���o<���ޏ��)Rpu����
�J�E����v�p�׫5/'q�D'�&I0~[ϯo]�5]v��j�RC&���2���ɦ�=�p׬�a1P�mM�hF�$ g]�������̆>����!��Q)9P>@L?<���m[PP�~C����֮(�(�H�}��[����V����C�Z�G�0���`�67e�;�������R#o�YC�?������!C~���Q�.I����,ު��;�d´�aO˯Cj޲�ө�h�٫G�.���M������ ��ls���1(`��QՌ�̑UUz���g����~CfHO~�R.��n��+����w�����׮^o0/S��X��a�m��c���$�cd���c�~�FB�G�t�s
�Q0���ʐE:&k��
���l�\�03�G��&��_���
���'�o�G�G�aX+&h���B��$4���5N�D��A��"F��}R�ϻ�T"̇8��=?a���j#�:!�b����M�6 �<K"\�_��i&�N���#����R�@� (]�d����+J��4[!�o��ѢB�N^�~�tZo����&m��A5���f�
h#\ްŹ��K3��<�t
��Y��	�<����E�na�n�#%�7�� ��!pKf��I�y0�~�i#�0Lu%=�%�
��#3E��;b6OI:�:�YF%_�����>��DSws�y��z{bl�i;�/*٠�&�W_�J�\�p[�=!�'�q¥1�&k�/�j���9${Ab�M��=��ߔ�>��q��uj��cF������s��:V�ht��z�1x8?�R�RA�b�I+�zbTP���IU�U��v� ՗�UJ>#������Kaf���Y��b��վ�=��YRH��,�,۬��ኁ�ԡ����I3F�&���f5�k�
��2=Eu����0GN�V9�~��DԶl"9ff��Y�HtJ���_C,��a�U��pZ.��p��M\A��������(t>��eތ�MkYo>� ���dt�\� ���]�.�SL�Z����4�a�(�*����^鷜�-�ٷI@�
�@�"˨D¥��#0�E����*,ƌ�'�t�!;�{��U�&���=�Cl�2�p�t4{����.���
���9V:��3΃IO���^C�1X�ygq�W�f/���qѥ��u��uq`^[b��şB�͔���,8�c��R������i[��瓸Y�g88iMB�E�"V���}�h!%��;�p'�В� ��<��;(E�������a�t<���(�k��i�NpFu�g�v>�A�În�Z�g�u�w^q�2��h�{��lNT�kО��p��Ţ��3�&������/�q�I��hz-���n�6�x�m�*ʳ�.�'���4#-�J����Z�E#b��l|s����q�|��Y��7f �be�y��#��E1d���=#n���@u66��}yX��,��J��}�fO)�环�w�I�_�6S��7�n���"\��կ�kAC���Vu�t�ك�C�}��R2v5V�Or��Ž,��y*Wj�D�ۗ��d��T��+�!4��c�  T��h��^��
�[po���Q9�����z�}���R ��I��N���zA%e8 zE��V�oEh`''Zy���Ep���(�Q034����H��P�6�k�X��*qT��m��<�xɾ/�!|Ĕ��B}Y��n8�z�E��n��g��� ���#�T�c����Kj�IFz��(������7=tv���P��w�������t���T�s/i��ն��EQSk��$�y�v�_���7�.N��/��|B[U���m��uX�=U�>���˾ILW��^ɤ�.ƽ �2T^]HnZ�C����V�bD0���9w���M�9����[fcF�:g��y��R���2��:�a�ps�Y�Z��2������h�d9P���M��㍡PI�IM�.��_��A$� o�:g�$b���#�S�X���8����ĳGD�X�"k!�G�WP�,?��8�Բx�^�9snN��t�0��h��~�ߣ����:ЄX�摟��`S���콎D�e�m�ov�C2�1������.� ��8��l-&j|�'f��Fw�>fȄ������фשBc7�9�L�`�~��WIG�>[p������xl����h]����w-�b#��n�r�w#���m��.���a�!s궁�1sN|	0��qw���n�Q�g7V�<���Go�`?�[�GM-��6y>W��?Ax��-Y�Nި� �c�c�����E�<�kB���$w2FwN���߆��:;�=Z%FD��-���F��V�	����A+~��Lgm����bt;�B�0��(8��[�'�oi���8n�4e�Ϧ�P�*j��s�8��M!$����LtBu/E𙂑j�_PAU��궊��vg l��ɡ~5�����O-7�,<^��<�w78���l+���F���	e꿳e2��I�;�sG7���~V�r�
��nG�X�,ܷ
��NQ�0��s�@�k��&}���尿�Ja',�3t� 8yẩa߆Qa"S�����܅Ի�&������/����+?t�k'l�;T��~Mw\��+����ϕg[s��(Q���%}M��L�d�@W@�����{'���o���Ju��[[��4e=F�8�"�P|(m�V�=�ƪw�Ob�ڀl9s-���;/�٩_(�`�*��xwK�]S���������=�R�qW�د3Q���[Gܪ�:�޵���!דm%>�/g�׊�_��T�@�n��4k �v�t�yڨ��bP���_�m#�����+Ed-�f~&��S�st���;���W^�Ֆ[���L��MUz�(��Qs�y�������S�ΰ�r������giA>vqk;���Y��A���{*V#d����4�:/Z��V�����7Sȣ�[�yr�����]+AG�諳)�m=� ���A�B��h �8��j�"=^�P+�9�r�C���F��e�q�U=��o�.nv�PJ�6:����t珛�W���)�6�r�~�[앶���|e
�PxQ�e�G	�hsA�Z-��J2��z.#�
�@=���M��-��\���9��8�)E����2�i�nw>@0{���n���r�����G9:$b.5���yT
�E�r�Js>8������H�oc�\�ݡwpZc����U)bh=�9��D�S�I��\0���P�3�YexvR�)E'�v�ʳq��q1���9��?Y@�8$Mo'���ҥ��w)S�|�#�q� }O��J�x֜%�s9HKa����}�1�@ԑ�!��t��6������[$j�:�p�C�˶;�`~ �'�[��rͼCBj���be��前����t�x�F���2�W"ă�y�T)���Ӌ}<����KD}S�yTf�H�LϤ�H撮���;
�i��J4`52�=��Y6�<ҿQDJ��/ͅcȩ ��'��$�^\����9�"U>�gzb�#��>����AA��C�[�����ȇ����O�сs{��[��>��]�#�#{%��a�=u�,���fs#v%�$��G=��Ã~�N�U��73e�a(���T_�hV��>�h!����$2����wR��q�Mm�8�ַ21^���Q;BO��;�4"��P�����M��k�I������q�]���(�P�y;�tҌ$�������QRp�{� �3(�Ƌ;�Ajg�&���֩&���d8�J͒t|kkȵ����y vzX�����mwi���\����C�^,S�0<��>�i>��2��Dhw*�}�.��ȏU|1��9O����1�u��Z��a�RAP��pS`��/����>"��Z�a}�[cJ����ݔI����@{%C|�=�a&�黈� ewPa1\���FʃZ�gX6��<��%҅IH���38�y<s�!�����X{���\ɧ��$,B���Z�	l�2�"�˕�ܡ�6*n��!�)ϣ��x�
���c�m)ݥ����x��n)�7tb�f[	��Ng�}��E�nb�_�P��Lh� �a�u�ku��n�jm�р�/]��X9Gr�r���Pgm���� S��f�H�X���'�=��t�Q�]�5��5�k�R�'��C�yyCޜ|��sô6��[m��B�J��,�'��[���ț�)�]ѽ�WQ�<$d�q�4\��]  2l�o�Hr�?�����}�׽�k���D��l\��1���K�}��O�R�?�[��}'Ś{m�-f�-Y�y�sA����S��5��|z�6�e��Xp�~\�^mf@m���퍧����T��(��e�>눶� �ۃ����(M��>����f����h��~����t�ȧ�l�&i�]�
Q3�=���]���a$��1I�-O��=�M%9�Fd{��5~�M���UÃk��t�&�Z���7��IҤ�@h��YC��<k1��BN��fmb)��9de՘��$o<{�}IK)Є�r��d�ly0N���Aƅ�KtO�Ƈ1B�X�d����f%�GD������uz���}���>#�y�N�]}��ng�e��jDK� �=MHv&��t�����LQ[j�讫��M��Db�~�M��4�l2a����qo�0vI�o�T�\u��<b>5���W��Jx�M/7C�ZD�Ťr�u�H(�O�~�b����:���I��[D-�)D]_\Q�f>#=�d.���N�ڎ)Oe³�/C�:���p���{���-�s5��F2Qk��S��u*�h�5f5r5�]��RIG%os�],�`-�R��0UG�%�5�mr�.���<UE�P/!b���ꅱ;ђ��<�* 	!v�zP!�,���F�%���RfH�>,��ڂ]	�Jz�4s�Oa@ȅȪ�6��kh���[�FU��ù���q�����!�)̬�{w��v�$��hG�</>�ֈn�1�������Z:�g%+�m��qgB������+t�_ K�΢�g$�m0J�ضԣ#SV�|�H[�\ȴ�£��<l�{�b�}�d�wk��3W�I�y&<ba�aV�Q'����0����؎�%��ƴ����_�~�z���S"���������}�c�F5�ˢ����0=G<k� uy�����HZ>�X)��CI�ϟŭ��,ӆ<kS���@X�g����ş��[�V�}'ܯa (\�V�R�ʹ�}�� M$Rd'����QD���oȰ��E��Z��F[r@��4����?L����y� X��d �*��+ݱ�T�m������T���<D���ѯ��ݪ�����Y����4��qv'ۥ�� ��z?�.�3V����
lpo��
�N��\Or����Zo,=oDĸ\)���>S��I"50��7���U���CD���a���{���U��㝹%}�5�7�n�E�X�� 7�|�^����	�Q

��ʩYƼ2�g����S�TA(�1�o	c�pVc)z}��a��0Z?S��#����d>��P�Vn� >�q^{��Lw�	��;O�B�C�0F��v���'H��g$��G�Y���T}r�M�0�޵�OK�'UȮ-s�?���OW��}�C�7����O�+��Z��UP-L��&��pY��'�(r�x�������k_�~�{����'dM�ː�D�2#0�"p��>���%�����wB�$��#+c���8 ivI�5�����aP�W&��NR�1Z�z�-�bΙ��Ce]��g��P[L{��Gͷ�f}O��w�,Ɩ}2���?��(Vm�i�\�#d��+�n6>}H>s/+�+L=�]������vХq��GE�-"�k��Qױ��fMH�x�x�8:~CU�  Z
��(����aj|��O0DX���-�1�����_xѿ�p��&lL�HBd�ÄA��i��uį()T��@Aō�1Q��b���KQS����pT48P uV@��oQY�[Xz��U`%,�S/�xi�fe5U�jvT� ��%jL޽���|
`哔z��q2c��T,��1����}8�se%�����s��h����>5�����6��"�(��@��Ѡ�W���G⼄ϻ�J[uPr��
��>R\�0P�a���׵��J���w
6j��cB�o2�dS0Y�?:�C��+����ѕu��%^���h~��{����x��$^��k���G��/���sQ��u�36�Ɠ��:chv�^P��o�o;�c���F�7�-}��jA�!$�L����(_��Nz�77��E�B����r����,&��I*�	�Kķ��!����D������r��;�ʄSIi�O�|����/+��7���hJ:��8S-�{e�Y�6�4��9&�'�N����"�񯞉o������n���f@����,��j$��L��4*��.�Bٴ���kM���6Ҙ�] ���ǒ�r��̄sTu��>9aݷGvd�!(��vٍL���S&P��m�B�-E�nKa�a��$��EQ�n��C�^Ys� T�<�� N��L�|B0�)��YZǲ�����T��%�f���U�	l�ίy#G3}�:`���ԕ2p���}�,D�'Ӯ��g�l�����5�>c���f@���K1f�Y3�!�T�:H�Ǚe���Y0>-0�T��1Nu�X�H
*q��?�#��\����1�B���o�C�C�]���>��Pr�{{�)m���1��^�yئ�¼K��@�]LpD>k�t��Ы�.�z���X�j*���o4�uؗ��dpӹs�}��i�D�O]����m��9�bvzl���Uu�����-��)�؆��%Ð�R�s�N5Q 1u n�����������i��ÜK.�ȇr�|)ĩ%7[��.���([�^�7�����3܏�w�(���wa�7�1<�t�+?rg�d�6�rx�$Qϯ��v�7C��iz'=�q�&���%E�������(rf������0��~�a�݄�#dT���ݲi��]�R��
�2����d�6$��%�eȿ%��+�1I�9iQ3ї�r��F<%&�Ӄ�6N, l,P�h����7�Q"����$��������7�+'��b-��e�YB:��\:/f�D�H�O|�U��Jg�S)���}&�I2#8]�eE��Ƌ%����c�{�nbG�
߮��U�=�F)o��Fyo��a竝�&�ש����t��LE��Ur`�R�|�j�J���*����K8���Q'�:�ò�,�Z�������J�O�
�+k|�%�/Lk�&ɚҒ*Ĉ��wmd��ۊB=k9^��=��} ��g[�>�̭-J������Yp��"z����{ZA`�A�+w�4�~tg����B�t�N��n�ǐ)�S_�wV�8�؈��z:����!"l`�<<A0+>L� %u�u�L����tږeL��MD� ���
W�Oϟ{u�-I��ju��1�(�B<@��Q�g�M�zż|�|	HK�#$�8gH��]�n����֨�DIiBBP��!�敜�f��z�\)~H�L.�N��7jt?��_���µ�_R��#o����+�	=��UjAJ�_��3;���%o��v�jx�H�/׊7�'< KؾrWC.�%���}��!�D�����'婈��f���H�����HqE:|}xQ ϱ�/�*J��ďy)S,���K��x�CdS�$|��q9�v�"���˄y+���U	x�Z?���#;3;WJ�R,�*v���~S w<㍸�y*��y�PЫ�_t}?���\ P�\�,��|��gf1�YG-�������4[C1n�v�P�3�oW�I�ҫ�^�9�e%��W���3�Y��Ɣ�	G��5�'L#R���su#��t���?(H��dV��p��l���!_:����=6ϩb	�� ĭӋ�
K ׯ�h��e�C�:2�h�3�1Z�d���>w��Q����J���{����(��s ֬�T���K�6`j#�!���v�"&n��b�h��btn!`?|3Hg�5#fz�;�.ǘ�c�n�h�nA+������T�oĴ�r �K:�9����ku.��3�\�JPѦ$��(+L  E�T�j�tV�Û��[I�]�D��$jtz�F+a�JF&�l�
x�/@��%_0��Cn=�\Q�Ը	Y�SDY�F�5ē�)Pg�^���w�9%�9ˑ����덣�o>DO�YS���<-�*[��s�-{����#��*%��������Fw�@���j��2�궫x߭���V�g�Obn!C9r9DLkh�+W���.�X�=�]��%�v�Z�L��A̶��(��B��+_�)s8.�{��-�铜��q��Q&�G�+�������`bz?j����Z#�j.��%萂+�o�|�Tfe@�����4�ʲ�!��DuA�.f�ܗ3!�C<���&he��Y�}B�`ѥ���R"o�Ɲ��1���������p+U���X� �wI�O��1��R%�ܵ`�@���T=|O`��c���"Ϥ������P��Bǈ�j��q��ܻ����F�Ē|�+�t�Gt/��QƼEP�qj�8�@�S%m!!��1���o#'����5�2����\�C�ƪH*s�H�X�����l��]�VI^���a�m÷��=$�e�����0+���"E�U���-�)	q����'G����MH���|
:rǒW@EZ��H_�?�oΓu47��F������i8�/|���� �#bm�:�'`����r���.aj����
��
�=G���ɡ��M��]m+��JgK��4R�b��e���ᕹ�N��N@�ǐg[�9P�#0��!��0![?f�;I8�C�S���p㖅"���>XN���R��㧑u.�߶p�T�!�!��\����{h�p��}2'�)�.0Г�x����d��՝�"vIVq{���D���I/i)i���,d�(�T�Tf{M�3�d�iԲ��A�lCĆ��.�*˝�n[�t,Дri�8�.n�}��[4���R���f��pݘ�ǔ���92&O�~��������J%O��Nʬ[���Y>Z�D��	�wc�`��Y��z*� HX�Y����8�{B��H�Ɔ��f�U�f� ^��=*Ȫ�g%*��A:I}C`5L��E����ں$�?/��BdI��b�=����6v�h�#Ss3�U���Åg��~!8,���S6�����ZDH��y:Dw� ��^����0��f9��Ӫ�$a��g:���ޞg��}�Y�Ƽ��3&<��uP�lQ#1p��
lCZfKL���})#D@ 3�=��� ��X��6d�:iW��z ��`}��͚�jh�q���[�3�����2$���ٸ��f(����_�K�
-L57��n�>m��g-M���ԗ�$j��p�%�BM1�E7藺~�O�ø��Y�\��U�Hh&�ܳ����_��� ���PS���TC_�g��|M��}�H�tqm��n�H���o�bp��l�VhC�J�m���95}*�T�rJ�kO��}�x<���'"ڞK�q�t ��uP�Kzu¹+�U���ڊ�����k^~m�:�1��y<���q*Mu)���Q({3СvY�{I-D�����������5�|���>?ƣ�o���� ���� C�������9C�Y5<�zY���/k-M�Ha7 ����W�4��\�M�l< >{��Kz\E߯�c�G5�s�zB�@�/��`�=b�k� Q����R�(�p:��Y̠E��[�zb�-�XV�'���-�<nؓ4k�����!��*Fv�حش�H8#�?ʣ;U�<��̐�g���x��1<�����RFm�z�a�[�*�<��K��8�}���Ye�h���fx�f67P�9d��{�b�b�/>d
��/����G͜���$���U���\>Z+l�70/k�H�CN�w&?-�܅�H_'�ɺ��S��Hc �9����pmcl�_�PʴЋ�&�se���l>��e�̻�t�a=��5�Ȃ��N��NW=	�P��jh���A��n�`Bt��Y����A���|v�J�U��}���l���<A�f��df�в+���;A�j4�;���m�]��rҷ�i]���d�K�Y�~EZ�uAқ�p��*�A弦�r%߽tj�V}R��D\�����ًp�6X\(y4h��B6�_ s��MV�3�c�9��!�R:�'r�cst|��,:BL+I+����H?�Yn��s�y3��@rh��)(��>zdl�e4K��X+	Ҫ��0D��i��{��%�ܽ��
i"�RF��O	�_հY�^'8��Q�����(����R�� �	6x>Lk��õK����z�$T�Tfv��$���l�#� �`U-+k�ρq�}�	p��mBKߩ��~�!T�tN9�\*��_��!͇�h�N⟀��V^	zI�q2Ď�A󽴏��H��nv��z�������ڟ�s��>P���6Tu�~����/�9�����u�����j��?Iu��r���W�����ﻟi��倫�z��H%�z?�t,�VE��[��t�� ���s9�_�M�DvMl�FnY X�w��0R�,�K���U0�B��qɦ���8:�����G}u�ETB�coL�u��j�Q�UT�����jն��k3��4��b�H���g��B(��o�%�w�-��܋��ܶ��S�@�r�x$���������DK���Ϻ�xێ�AW�M^-�������c��|ߚxo]�v���e�a-��\�}r��d�$���?��b�o�Q����a��\F�8��>��A���.�����Ƹ͜�� ��OC;u�D=zF�j�H�^|� �|��%v��ݖ"�AR� �X�m����#\k�M��Y)�r���h���К���@A��ޮ���7_x����]�G�;מ�����;av�EIc����*N�rt�������__�S�|�v��93䌩�Q�I�O�q���v#�@9�/Pfz�M\�L~vD���P� ���g9�V�k��%�l�[���_H�-{��lc�'X�7B�q�y���a��ƍ��Ny\]�&�A�!�s̓����?u�.�$��0����V`'e�%�jx\G�*~suRY���g��Y��Ȯ>Oj�����4�ؒ��`8t��Q4)U%��r%�S�M����JcQ9y?%^%`��JT�6�4?�Ɛ�I�`���:)/JB�}	��)tҚ�@��+#��r�뀫�,J���wʍt�^4�4�����[���b/quh��>�t��;�w�a��*�`7�9�����ɹ���p��g��9sf���|S��c-dg%�N��N�gC��v)P��O�\��F�m�#){��㛜����4^�"���9V���6B�-�}mv}Z�(�'��a��Y:j�kԧ�����~�Q�hN�=EK�(UVHG�i�5zv>߱
��m�6]��+�ڿ�&�N,��i	2�;3���O�"��.�*�FЧ��c���A���vA���:��ϙ�W�us��B��*��zIO�f/}��<i"�"%|���\�ڇ{��	G$Լ��d�uj�[�(L�?iN�OW��ŪR?��>�k$����~2S��V�Xp7�����]?L6�ư��p�"[:��������s�eӒ��Z��`0���{=�	���wk�b�����#�1�P�d�n��˕��&�H��0�@Dvv�U�Gu�`���LD)=m4�F�c�E�lf���  �q)�7n��H�2{���S��.�C������oZԋ����3gσm��>���nnkN8����~���|�ʌ5�ϼ�,�C�Wo�Պ�qY5*l���p7��/]���7O����?BG���.l��l�՜{F�� ^����Zm{��H力��ysۧ6PJ(W�#����7u����"��TR����/���-�����Q�{m�8���C�ߕ�R�Ó�%�L��@M���Ȑ�>�p��q^�����I@�82[�
A���3�Ż���@��z��0��"��|�8?��y���O��×)���e�8�ڦ����C��
H���!]�p���F:�3�eM��y,r��?x�l�}��tI��>X�����:WM�>�`�÷)�=Dg�&�m�Rz׃�[�wƤم���J�p*��p~DMҘ4?y��̜G /��L�g�s<�E,^�Ð��
�F��
X�$��Ku%q/���Q�%]:����/���V��i;���MX����6�;<��v*a:<t�.i�. GT jAo���	d؞��f�Ndr�UDR�:c��u�	0���t���aF*��m2U��|8J��{�"���J�U.���ı�T�"�sM�cVe�J#ǣ��cgj���u�t��=r�t�a��m������	`��������lvs;7t諈��E�ݧ�Ps�)xU����X����e�XMU�
�ȉצs�B�Y��l'>���<��{��RY�3�4��<���Ih���4g�;�)kq )�U���Z-�TYW6����F�' �?m��a�Ӱ��/���Z^���5�y�`O�Վmc:`�Pr@(��ea�ǻ2!Ȝ-1�+����{_�=��K��{�9�2J\��A ��݂a7DP���}JO���0�hzޕt�ʧ��o!�lpyT�Ft���{w���b�`��-�]y7f��N�Ep{������rV�)D�w�
��z.���dzا�Z ���Kū�, �����|��$Ɨ2�m9-z�_�m��<3�a]�b'��	��͊�H2�:���Z��~�y���m�`*?:Xav��U5�$Uں�d����%������oT4c{D��ь�Wov�*%R�}O�$����ge#�@�r��n�=.��T�v�b��� Q��
��?�q;W�W�����g�l|#̜���>f�?XSN�ۭ�/���waLN��ejR�i��u�A�J+�{��o�I��Ď7��	"(����N�/��Tz��q�E[`78/O����vU��xB}��}����y�M
P���0���:��jJ4����x���/4XYM��
DDXR%��it߼�^��3�s�a̮��Y�M4E7�\�P �	�ik�)��l�7�b�s$��Pp�zT�j]�+j�����˞y�����@S[�Y���٧���h��Q[��Z?�Eم{9�.DV�u��$�/�C!H�ټ:���$(|�OD�r���^�xqvY��g�����Q��E�
9�� [�!���$,��56�8ݙu�+պ����{&%.T>�a~zy�+} 7}�	up8;!ݯ;{��^ ���T��J��s��_N��zc�К[�5�S���$w��f6}=���h��{�_��'cuØKj\�{�ԃ�Z�vV�ؒ��Td�x�]�I�ċ�tɁp��q)�,�]�2�L��L���n(�u�����<.g�~�`T%�AE҇ʚ�J���^Hҟ���29|x��	@�Ƿ~K.C4�:���L��jD���Nd�}��~t��:�sU�,���{���S�Y���[}�YY��{|x~@�7Љ��|.�'��y,�ۓ=��y@L����Ñ@�k�D�I�˭ ���-@��*w �X�M͎����z��1������̐��EW�*��=���ګ�:��X� ݻ�ޥ]�xY���>۟�2��޿B+�&S��K�%�=+��u�)�8w� w�5��F��I�r�B���W'Ew[��ʖ��Ѕ!�����R���]"�kԔ��<�!{�^�9�ل��g�t��mD_����u��c��҄�*'+�e�O_[�cm��I����	62)U�8�=���e-g�E���pc�m��t��49�čB#<Dn8� h�O{PQ.�ϡ��ʳ����J�#���fA��8��Ż��q�4z�Pi�M�86n@�'LuQ�@Vd:�T��4	.OhɠA|��4D��ٹ��X������;)P���L%F�JLEڇ����M��j�O�/�i��8K�Ҋ��љ��*��62����2�Ok��X�&��t�¾ʆ�"�TJ��/���Y��Q	�K-��O�$��NF�p�a�*Z�T:|j��gciD�kdG�Qa�T�@o+y��yG�s:���lU-8��z���R�7��DU�]����Q	�Bl .���������C� t��`!lf�x� Uk����aV�e�����UP.n�G�o� 3<�n�&}6�9�r��	�A��R���k�D½�a]˰h�x�CA�t|.�N���D�h�]3(][W���j����lY[���U�����P<�w�@\e76���<�}���g{�Su��è�=z4	��;|τ��7D���--[�,� �_�����D�Ng>:;؁t���e�W>:�S�̻�zpr��Y��(%G,���^�j�s7/�����4*��̬�؀�b�L'�C�}�5j�X^��u��[Ų�P��NLc*�0AB�B��լ|�R�T����]׬������Ɓ�`�n���ե��\X!����]�_�x]��\I�}XY˛���B!\��<�F�����E���+P�Z4C�C8}C��8fkG}�5$��j�5撞�7��JspS���S/�ǱtQ|%\���{��s	�@�4�|��%���e,̰�Ÿat4����.U#����CZ�����Ie>~IQ`����N\AB<���9Y���#�}~{�)k)�����f_��7��gx�H,��!eT�Q��	�	l
�y���`�����oas[��CT�z�/�z@GD�GQ���:N5N��"��L� �v��?&� �-���Q��}J^t��n�8���x�
�ɓh�ad�r
}�J�`QǶ]���/��f�L��o���^{�q�Ŋ�Mt�Y}r
V%Q�'�?	�&�QY�Y��P��a�;���>gz:'C*LQ;:<��=|�i�_[��ޑR)l[%�O&,������A����h\�ڂt�g�7�Tg&�W�؞�9H���{�h���k���>�:��;�Fc��F?Y���w��zV�+|��ˆY�E�1'�}�9.5����\m���@O�^���N��ہӞ�wi��8���e1nv�rĂ�����n-g�3۔��ԣ2!DNy��1�խ c�3ɕ%��ݷ��T��+ͥE��Aw��1�	�l��Y�P�k�\qzŦ�xO�P{_"Fڪ��Jn�K�}���X�2a8���]X[�J[��O�~j����Z)�#��?;f��*Vne����:�����28�s������_�C[���Q3;�nmVT�C뾣�/+��Uaw�(*ҁ�~�j��ְ���[J�R�I9<��;�K��,)b0i����;6@K[]�{A��B�<� ��rYb��N<��G�j�|�'��������іCN��q�:��׻A���d���bn�ճ>���w&��6�����R�]ꍘ��צ�T�:��ӎ��hPK�,�|:e�������&:Աt��E	ˎہ�;>��͠A�'�F�S5�X}_+b[�9��1O�!�ʬ�F��}G�@ `��XU�{Yf�\*!t�nK����E�q[����?�Ҫ�u	l������F�h9#݌��d��Y)}Mk@`�벣d�s�����P�h�h`�i�	\��8����Vٚ�h��ݻ��t@p;�տ_;?����`��8r��G�(��ޫqZ��67����r 9:"��I@�0�L���&Y����8�Aٮ��6�
s�ڏg��c�ơ �����}gK���_ ��b�ZK��p��r�t�ׯ�����H�.3W
.��?e�<�3�6��0�'��N9*(�<���)� }�ހtF)�#6~�tbǽ��)���\̢��J0�>�b>-=���X��Dޔ�!>$�U$�/��_w�Z���Ay��cGZ�m�AF�Ղ�؎�@C��ۊ��06B�-r��kt���(H�];�d%���J�R�M���:^�?�mI�/�Ew����|G��3��8k}��oO�Gܷt&��&ŜEJ�U$���idB��3���`�c��T(��8�*AN����!��zA���|��~�$�cY둝x�Ӵ�B#ñy����`�R�1���>����M}��A��S�K�\5u�L)]�eci�z�9}�R���%OJP��TE c�a�����lkgy�Z<Μ�3�n$�+ͷj���O��l��Ұ`y\��jz�i�ʵ��6��@�ж�{il|�88�B�������#��i�7}����"!�'4�c�}�A� $��N����KF�T=oKr������$Z�N}O�T`��d�gClÀ��N�{���=�4jk'��R�G,}A������3�Ɩ7(.�K�hU��i��G[#K���Z�}���Rl�Dl79s�s=���ҤcP�����[�$��_��"_��h�߹�U�������N���TL�,s+]O[]��v�yd�3�v���Y���%Mc.�g}���n����Y��jBD��,^"T�5Z�qU�U[){�a�$ME|��^A|*�|��߾��i;DU!�2�ɳ�S+�{�lQREe�s72�}�(�+ݓ�s���#s^6p�����6����O�g`� �`
x�f��0}C����ߩ=+���%�����G&��ៗPj��ˢ���E��W֙�lu�d���)�*f�܄v���$�|� M��X>�;A��cO�ldɪT8������-���|��&v���Iv���V[��2iO�`>^Ytޱ�-g���d�'��L�ݛƣ�&���k�8a�(��+�[O;N��^x_���Yٜ$�n��uLKSd��.��|[%t*�b+�t�����������Ɩ����x��1���]ߣ]��q�f>��[U$;|`�\�Z�F����M��`{+���@����E�O��݄N@�#f2�ң��1��y�;& ^.*��_��(�5����bR&KP��@��k�n����{^f�������g���0��6FL�J�_�������ޞj��X=He��5���|V�{�S���1dKa�:�3��*L�J#k/h�ψu�6|D��I�n	�JC��R'�߳G>���!w+��׶�R}��&�i)��ꃏV�C����VH����Ơ���R��}��|1����lI�r��,8+/e� ��,��0jW���;}.7�1�:��r	�Y�J@�A���ORc�t���M`z�$�t`��T�q�ǅêL� ��B�ݬ;0P +����`��⇃g�_��C��SP8��yV��-��^Lln*��'�c�����X*Ъe�D��F��lEoQ�u�-N��/S����9�r�
K;�+A0D��S�v�����H��ޫf��G�O���}�w��L�b�!(}V�*��'*��=��R.R��)��+�JtJD�J�<�����-}Q���0W���σ@�f�Y�e�ÊMmdS�;���!����݆&�)�e��IW߄�u��[�D�9����nq�pE0�C��W���#��P���0�kc,�)�J	�Y\U۝b�����"h�� p��1�"�'Te<-���N_��#�l�F:���!�cfw��"ܣt����)&�	r��u�ռ���q}!_�)GI���H����l�{���o���{7Q4�R��M�9�e�<ti!�,�'�Y~��X�A�x�Y�G��ak��}Qmܙ&y"^�����;�񧷀��~����hj���̛�.	f]OԴɅ��> J�k����}���ThN8_�r���n���oI�I19B9�*D[��W��,5~0�fZVG*df���Ϣ��֋#���!"{1?�{���@<I�v2���G�A*�^U����1��Ň IClw�4�%�r���m>m�## ���e����!)O4�ȣ��F��)���w�7�߆�C�^��>�Y���PZe����`�{�uPb#%��/�gY,��ps82�7�������|���7��\���l�y֘�f����b��2��wؖ�p��}n�4*����5��-�f< �v���$_��\##��:�z��4&�o�;?ϰ4�Fļ9��M�-}�c��^[B�"0$�3�$�ub�H,`R�|��Ϗ(�r����r�U��Y�&L��$�񍠁�����~�J�������!�|;"8M����?\���9 d.VL�ɵ	e]£�����P���A6\�\˵�����~hhv�.�x��Y�D��+@�S=�@�x/����7�{����!��8Ϡ�m-������ ul�s/�O��$~Nk��O���+��75��P(���~ܞ�� ��맹�h��O"�����M�aU5Ƕ��X:������-�OT�[,N ������K �R|R�|�Y d�,�+E�����<�Qǎ/��ԉDYf�`5(v�������Ih� ���|T����8K��W�]�����؍��p��|-������NxS��f�W��o����܀�F�y�1�}�5*�G7��Rѽ%�b�An�[z;D����*l��\���4�WZ4�"3s�+b��śE]��o��!N�������6P}�x�"�7V	� ���X�u���T���i��x�6��J��pLw~�����X�,�y�Y�#�W�x3��	�7�5�8�T)���vdI��()��}��Xd���}�q�ywY�*ƌ�3�D�Ԭ�"�H������m)�HueQ�&�#�˂d^��, ��_�y'�E�c;@B���c�]��ׅ+ 3-"���n�J}��?�z�ڀ���U��o%���%f��4,k�b������A���a?�#�)�Ÿ�=�`�b��j-�?lE@�m�`T�xu�C*F9��k6����ڭ�S	�sw��ʓ.]��[�A�5T���)�]2U(�"�p�8����g-~�#:�u� ܛ�T��鮹%�}N�*����P<%[�Y#��I�Ϋ��eυi�Ad-(W\��~���,:S�#����w$��H:�¡��u�@�q��c��41I����OR��3�3!)ٳ�(L.�tXVr�Őf˧�2�<2�f��8\��e�yo�^����= �ƏPI%
��fʕ�v�T{�r��ʣK�<�''ԏ���pV3_d���!@���J7��H`<&�ʐ�@�g�h���=��VP#7)1�P�K�A �X��)��~�#��c@���q��B�uzK�	�"=m��?�D�B��i����u�{8�3����y!�5t���C4^i+���z7�/=�69���jAS�ߌA�w*�l���+�@��m��(U��&�� �f�Ye�EZ��fɗѧ�'��'p2Ř�� �����Z�]���Y�FF��r�/����URq�
�9º1F��L�P��[�t����X��b7�F�N��lK�!4!�4���"t���ON�b#)�<��0�D��p���O���E�	%+=<��>h+�D���a��CN�Jx(�^�kJ��a�q���<���u'���P�zk�
v~�fp�7U��E����qN��D�ݱ䊞��(t-���>�*fχ�P�~}p����xa�x�L�Y�2�p�2kL�2��� �:`T��;n�"Q�q��rJ,��rS�}�Y�!t��4<E��8I��ҝG�P��;V.�]~F���$��<�sm��x��񶌧v���F�1�!��H����@��$4�5L^�����w9<��)R����ɉ�Lq�Qwܔ[ߩ�m����u9��FN)[�,g��!H�~�QNd|$ݙ2�!]<K1ƿ-�WG�k��и'�
-Y����"��D�$�����V	E��e�M~���J*|�
�;)z5��ak>F���@WP�p�	٬�p|����'j�ig6���%ˑ����uQO���΅���Q6t�-�֖����n�@���e�^��\�>8Km�����h��7�#�#��_ԣ�l���By��G��`@.���F s�I/	k�6��ֱ_��$�f9��u���W=�x�[�S��a����/[A�k��ܛ=�E�v�3�
!>Ý{���B�0�|�$]L"�@����(���>��S���(���x��h1c��d��!�F�N�&��r��y�"T�0�	e��Bŀ��7+95+d���e:�g�!�|,�/Z7��H V3���gl��*�q������"�f����Jd|��&����{�a4u�V:�*&���.�?���XS�,=` �q?�S��'��:E[��!ȴ|����ִ�LY
K���-D��w*8�jڕ���O�H��zE˗})�\���9�8��?�R%X�B!0⍐RJ/�����#c� l�D�UϞ�c�T���BS�KQ��y�<�(v'~���oЎ󴜠�r>���D>�{�+9?�����.T�.�ȝ������[K�Ar����H�ɏ�aA@ǽ眂T���$�S
���D�'1�@��'���&��֒R��̋��H.���B�Bk�������%u�Es����#��L	��/����H]�[ɼ�C���EyX�&5���
�z�g��w��?�|�\�z���	���%����#�d$s/km$��e�k���c���Қ�~ɚܐ8�$���'J2��߯R@�R���	`ee��h�RA��O����b���[��TQ`J#��l�|n�ix�I�e�μ�i�]Ү�B|N?��L�b3��f��մG%_]�h�6��f�ߚ�����D�	I��<@���2�	]��4����3:v�Hߏ����a֦mL�����
�c�'{ft{�e�9�*Q-�D6��A�_.C���A�;����(Y�זjڃ�H#�R�'�˜�D�4{�� �j�.���s�\A�Sǭ���Z��M�7�+��˲��}~F� R*k9��Yv����+��^	;�u��;�
.?���/O�Y����������9�~�l��;i;��,%�����$_�vw�2�74�P>�`5�9�gY��>.ț?����S �1c0���x��mb'�t�1��{#����cj�]�@;j@�&���$�_��P^cr�'�f�vG!PO���8�K
-F�5��Ԓs�*���a�(y�Q	ZƔ�.�$�X�8@�M��py��I���"�:�3��&�E���E�*{��O�G|�M"*�{�s���>�*���ԗ���1�Χ���~��~�ٓ[�/.���j_	63���/���m��l6��TCy:�1�_�{v��ZBu͞�7��ϔ���Q�!���Dc�V5�n8Z^�^��*Nu�w��l�֥<t����f-�SA'��H��H	foN[�y"U�Sn���`�W� !ٜ�I&�:o��z�R��c8%�*�o��:6(�C��#��7c	�ʪK�К!|�ԁ1��mR�h����@m}2ØQ۷��k��o#u
��y������f�Z,8���
J�u��"��Ş۠½�N>��XP��S!�?T*�N�Q�%��F��^S��T3��išL�sƩ6�S�B�PN#�_�=��@�<�o�t�H)cY��@n��~)~ ̗*�ao�{�j� �+�7�����f�|s�TED�zE�WW�-�8nU^��z�,zN��/P˯v�`:�ȋ�aOn�ɯ��2P9�7��4�y�e�ش���P���{��>;V;�->B�����ʒ�6� c����O�{��T���lPǭ��+1��h�<�o�U��V<A9C34WR���v��J�8�i�� ����R�Ę�a�?-�镁���r3������TN�	�ξ�x(�E����_�Rr�Y�I�����^GMUV�� �����0a�Ņ��0w>j��+�s���3�5�*ø��m��w�猝X�z�`|��MOi��y�l���@������I�)�Y�ܕ�({�t�ۊ����	�!�U��*b�b��[���$�����?{��윙��P�����'�tk|� ���"7�-�t��^zC1�k�Q�z�����
�`����gD=�$f���ރ%�q��)/��*�Ra��eY���⺗[q����K�>E��e��Ixs�͚~������A�8q�}�pOc�⥻-�~
hNh��~�$[���#ehɣ��{��\�q�#hB(�*��X�r<��K����<=>N�w X�6��؈dUpc�5���*��wdY�U��b5zը=@w��60�-M����EWP8a�ߣL�`�i�F���E�\��f'e�V���S��>�L�Ͳ���H��3�9���n���|�Pf�L�����ke(q�����8�mǳ��Do�O0oo97��HI�fVC�V��7�E8���_N�7(��['J��6�y�#U�a�1D��g���Ĺ���\�Nו ���i������P!�F��?�s���/��]�@�:=�2Vl#����Z1�R�Z5��~Z�b��}FR��&��"� 3��Hze�<�M�����И�}����N`HK�`}/-��eS��a��HZ$��X�sͽ��.9� ��N���c����� ��i߲�
9�(�Q����0
�y�S@���m{{�
l^9��M���{'�
PV�����'��?|��̭�])߁h��.�u���p&���T�w ,��HCrQ�X�<vq �fAD�����M��xMu�|&����!�dl�b���jثox���{U���Mm�0Č����/VO�-1Jg��w�A��>^0��?�}���w��r<x�㫥�i����bE2q]|���>"��@�WxI����wauv<7��F>��޾��Zj��J�e~G7m�o!�.���y����&�Y��Ɵ9�D���'���R8����w���_o%y����3�2��t��9#��r�g��3Z������PH�a۴CЀ~ ����
�yo$���X�˶�Gp�d;躋���5�]���<k;R��C{i!6�o0�i��W��[��)XmX�j{9�t��'����|�s�"�ٿj�5�!g�8cqx��t�ejf@@��6$���Y��tJ6H�93@���%�����W�i6����UCz�;A�����z�¹T(ܾ{��D�	=��Qo�JbdY��Q�l�g��T0Nb�/F]�Ô�<va�����U�wM�d�L��R�/�ԃ˦t�y���Ac�t�����<}漎�����П����v4��fV�o5!��UB��C��?��,�"Z H(u:��,��T���8����B'�F�u�q|�1�+���������CO�� �<��^;��&�jQcm�
I?�w��\)�	@��뢑a}��jy�셀�)���6S����4u�|���+f�]�gMM�{r�-K���P��4���VI�����.�@��.�S�$�c�3H�q|�C#Q�)ݰ%�y�=��m�}j $�Z[R|�XZr{����nfУ/�%�`i��~��!pkbD�N��V����(&<-� ���;kt6���f�CP�TۨC8!;��iP�Ğ<N�&i����d��[Xθr���E���ωD�9��Ș6�I
h]$mȳҒ�׹�}����=	6W���X�Ɨ2�M�W|�amLV��?�bI�˝ˬ������W��_DU*)8��ڣ$a�����
�_����c=�tVIF���*z�{��Ӟ��2ȱ�^�� ���<(;�S6�9�u���n*x��Ii)�G����>7z���T,HW�#Z:�O�ήS\rwɐ��B�2��N}e�8��7�¿�c5JZM� �|6f���L(�Z,��K�e��h����f� c0�d6���vﰕt4�u4O��i�o��[<��׻U��,�����Ο@�ʒgʢBy����6<$%�Z�@)��!@Y���,`Qt�)��kv��m�B��\NG{4'{c�ɔ�0��������D��Y�We��c3��KM���f�3�����J	�����rѬ�+�Ik@}���p�<�i��J���|�I[)����B�
��%�Ӝg���a��^-f�g�2��.��~Ņ�]M�N��<�m��1�#f�il Z��S��%|�k��?](�3�f�|K����m���>���}�
����ɥ��6t��N�T���n�
���g�5�f�N��{	��=�̄�ޞ�L6@����7h%��p]!N:�Xx}4���o�'d-�5�k��f�a.�pk����efH�t�6�]{K�Z��J��{a����(�ç��`���jD�Z�W���˅B�G3sӮK�3���B�}'(Ν)/�u.y�Ƨ��e�Cs���'PEsy�%&
cx64ZZI"�d�zC>���6��|�g̛;c�tb�M����L�����������"�dJ�10�-�G��5���ʚ1�z���f ���*����:J�ǆ�1�܁Cы ��(�@H1�1ы{�=<�y<�w+g&RČ��^�kB�%`�됰��	?T�L����wN�y��2�ǫ+ZD��-ܣ�M)j���y��+�E��`���M�ʥ�2�$���:�
��
�E�;�qC>	ar� G5��?��r�9aD�X�����X{xI�$B�*����bp\w7�H[�ٝ�jD^�z6O�MlB/�tj^�3�:%)��y�m���)�HߌD�s�����茤���<��"f���5+��l-3�I�N���V:���`�`I��B�0'��#�%r�	{
����Н	�NՙvP��۲�d�ܺ@�E�	_���ʌ�S��!H���Z�]��=&�7FW>��t�z͗���W�좴	��Ȟ^h�Gg1/X.�R�uN��d֖N970�?��y��s��nP?kbJ�+��H$ �ӷ��,r�g�L�3��
	�>_ZS��~G�q�P軲B���l��,��*��$@?��AX�.yS�F���m��k7�Mz��OxA�n�;2����eQ�����;*��9OS��S��$�h�e��{���p1TТyU0^C�*;�!Y��xd�\X�~�z�-�XM����Ih����Y
9H�F�~Od�ߑP!L�̞�j[����w�������$!�߉F/���p3��f����[=�V$��ý$�i���ц��d�ҰNY��tl��RhwSC��j�Y�[ަ�Tzdj��[��C�PO��H�Ĵ/D)s��X����/� �M�ɔd$��{��?7OSn�x�Q�C�t��F�N� 7�P�����JPgS��rӝ?B7���H��J��>F4�Հ&��G�<lÙ����%��d�>���_��͓����n��Wk�N{"���~�^����mzƻ�-}y�]z�Ȃ�iZk붞��$� �,�N�����C ,����s|�P�� h����`4���-ͭx�A$�$�fT������t֩A���J�"H�o-��^���oI1���[���c�Q!FEb%
�1]�	9��̧�
�U�E_F�Ax�π�ļ���d�G��̚��v ��o�2��q��BE���D
�޼�h�&�_qb�5��B22��ۤ�%��%J�|;���+J�`0�
`E�Z��+�f�t�����R?�λ���MM�m����іvǬ�`C��R�k�<U�d(tЉ\~r��;�ofo,i��r�ߡ�
Þ:�B+�s���M ���C�`�8�)P�VQ�a��;>^�j1�2woU�|��� t��l��g�V7��g"�v������$��ꄬM�wpSo3b�)W3�� -خ��5}�ȉ�96��W�3��|�GH�t�ھ�)�+ �Ьܿº���}_�VU���Q@��池��k�8���,;�[kU�-�3�Z��ԄtSA;���z�z<X�fd���V��]�*��SO�2��NM��]]����8WDI;���t���N�m�6Q�v!��>	�+���lHl�6�����YoAL0o��43��h�%{����'tw�Ѯ���a?%q��^�9Ù��|ᥘ��o�
(�^�~LՐ]�}��>gl�T��:]�{
�#!�q@�=��h�~}ӆ47
HL=��`Cʁ9tZ��Kf ��ʑ��I��U��j�o�N��tQ�1��u<�F��9�K1��f<?o`x�J��(�*���$��3�.�}ֲ�%��l�P����g�Y������s�:�XS���
�\\��C6��
���6�C�Ch�cly4�"� VZYۦ�f�f�l���za�
&/���h����&�8��%jI�=:Ĉ�e'0�t��͟۵2�k ����{��y���!N$�ǝ��Ib�90`|T�^Bk��&��w�p��ӫY�ٔ��P���8o�D0�t���n���X���9]�R���h�wO�����K 2�(,{��3�gך�%C��Q�Y��7ܑ �Q	c��x�M��¶s�+�)FrÏ2Ѫ��9`�7��8@fE�a~h�^>���	�/_��^9ɔE��-������9�D�[�G�ML�jK	����e�ôBh�!���v\�*�&��ؒ��@�ZxϽ/ǻ�$�e��rm�N������fbս��
t�_���`��'�ʈX��Ч� s�;j�D���r����u4Šj���!���X���9{��vG���i��d��fQk/�7�z��L�����(�
�5\�C2���d}��@;q5e�>o�\�a��=J¹�A���FD����]����FnS�&�����H���Z�U�<���_pk�ʈ[���3���Lxp8/��e�#��l5�L�.
�fk$�O�mm�6q��G����C/��c5	�g\�M\}vʟ&��!���0��m���kb��/�G���tVI��Ü+2� ��S�m��!A(���mK�f��D�Ük~�����
�ɦ��h���b=�"�-	�_�JF26ת��6VU1&��3V]$5���fa�(�H��Q;C�9s6~
�p_��,�^��L���%�z���ս��u���$�}L�/Ju��|u1~�acL��a
�w0N ���
����̾=`��qݩn��vӀ���SO�2�� yJ���zFD����sT�j!�f�i��)��X7%�[_�'�\W���=:�4gdM�c~<7�9��L�m���f�PV\5!~�OHu�w���"&y.�7q�	ȳ�Ic�&>�wO8BGһ��0�l�g�cX�Vc:�cI/�_/�s�td���+�b�C�2�����QO���#��������m%f�0t��.�0����� x��@@/Oq������+]���p
aM�fc=��H�U�8��{�!�a��ǵ�C8�o����0Mb�;��o�^]�V ��`�/���U �z0� )�;���]��f�0M���������M���K"�4&`(P"�.!}?�PNvd;�� ���QN�uH�?�N��\2W�w�_(�@D��j�s�,w�u�˙8�tZ�ta��h)(uO�E��?-�n �H�K����b�t~�� e@�C�j�H !�MG��-���� �C�8E����%�l�c�G��p��.Vd�z�S*Oaa $�`��a|b췢e���մ�i^*�P�BĤ;Z�hL�zI�h�΄^�;�s��!��\��_Rs-� �Y��LK_�VX�$��?��]܉=�2��l���֑wܓ������CEs�9�!�:�K��Ӧ��u�^
N��!Oy���{)>��R�b�]���+N�&��I���AZ/��	�S�p��,B)��
0�@�E°��2N6	`�@vK��gcʼ�֙����"��˙S޹�	p�����r;�Ϛ�E#E#B#b��ܒ|�+s=i���n�1�]��Ӄ�:��o0�\��R����u��;�%{6"�tL�'��D����qF�=�+p�}����[�s�o�����@�"T�2M��C��!�͏��n�4�yD6�E"v�P�3G��p�&@����% �u�e���I�T��EB.��щP��;����DJ����$ո/�FxE\���j �ŊQ��X���QV��C~�C��I�&����13<�m~�Q�>U�Oᒰ̍m��S��R�'3>#��P�?U�Q[f,m���`#����*����\�����.lwK�;�1�V�[k�K!G�Ǧd+-��颐u�:nPp9q����<�f�G���FI���O3Cn��R"�;kpx�$��c�G��8��:ǌ������w�xM�@�U�IO�G8�ҦJu`��i��^#�'<���]���]���Q�Δ�r-��̝��~�ͨFE�$ӏ|����T�e�&Z���m�z-�����NM{S&!
k����®M��}M�'�����7��z��m&F�8��)�˳�||E�>�x?�^g 6i�`�^��5B3�X�fn���[�ƌes�Ӡ�ӡ`=������������H���:��� �͒�<S�n�d3����Qӵ���q����X�+�q�E����=p�l���毚��DQ:�-�(�ߌ;��OX�*F��L����8tOS��ˇ�B�#�krEI*�x�Q�Σb�v��>���8qb�1UyM��P�,��=��0^[��'d��`p�,Q��M�N�ɠ���oB2?bOi1�9��FF��/�E1+\A��%��\�n�� o�q�bCy�h]��ͨ�
���M׍5���O��{�1��?6�<��z�΃$e�0Ȍ��L,&�}���k�p�g��9쪁6~�/�P!/��:���b�e|���t�'��*cR�����:��3��Q�i孧�2�y����RWL�M��Ԫh�N����^�@����r�p#oq���͝�d+x����T�aۈK
�GK-f�~�q�s-،3!Y�q�pԲ6]�l���U�5�6Y���MG�U�[p�P����hO����1_�6�f!=��`���&	�Q�"n���٬B�Ϝ�\}�*�+X��Y#$$v��IH���-%�줹x�V�*k��@�0���t��G��d��a2�1^�ꞁC� ���� p���~���.�d����ɗ}��Cz.���Urg]�V[���C.��^?QN���5M����A�,��%@�o�(����i�\w��m�s)^�'�\��LK���S�ѷ��u�'J� ���xk�2��|̠��=�n,�L���p/�猪[),����U�sc e ������))�^F����H��bz����G� �(D�tDa"�O���QtV��@��oq�Q��7@�����¤�ߥ^�0azt��AR��;�kpގ{$��l9
D�uu�J��1'N�ʼ't=��qS���{%Fb�[�t�����<E���R�B6�֑?X��|�/�;��R<VP³����j�/|7�=U�E�)W��?i�N�0�xw#���?i�y�>|r.j�.�Q�If�sj��G��C!�(�^V	X]��~Ҵ��K����5������ș��(\4��Ўd��h�	>?�|�)ڳ�蛛�E��t��=�͐y�:HS/�EH�Q�ʱA�z��,�������������`Y3�����|M�Z$'~E"׽خ����F�4+!O�a�}DH a�t{%6�z���9���. �%5�;�B����"ޛ�4O!�B���s�S�$b�%��-0���7t�ھ#\��+���eS����{ �r��L	��O[�>%(���|��4IgWUNaOlU��o����+�p��qA���ܢ�^�9n��&�,�G�QX�<][J���:*��c�8����b��ħ���Kέ[�'}��
s2X[�OvM�F���p�[x,�����z[�OA��W�R�5N�##�KJ(�	�Scg�e*X���z.'?��X1L���ա� ���8�2�y�|��ǭ��G��Ai�o�u���ѻm��S?~�&WTCl���^�u�o�z�k��)��P8
Np���!Ɗl��Z�������HT���@�L��AͿ%T��L8lF7���V���ƟߊHx�B��=aN9_�_��|=Z]m@g���*����Do�{Sš�VzFI���Io+�h�;�%�����x_�5���6���|"Ė#C�Bo��)9ƈ�p�!�P��3�t7	���KW|M��Z�m��-G�^J��F`�UR��t����+kd����P��p�Z:��3ٿ沃<��f�n�*,B�(��$�������j���Ѫi` �:/�P��.℻D�)%�v��-�kT���M�mc�CQ3
k���ץ<%_x4̓9@j<���h*��������<o�����`���{	s!�x��M)3�0��C�)h�a��D��A�]�/D \p�Z7u�s%�OM��dz�;LJ��g$?��c;9V�AjA�2��M�����,A���},�V�S�[7�7`y�9�Qsc^�d2aY�i�S�������r\�(^�YwЉ��{�y!�^��3�H� C|�W ��۾f���{�K�E׻�#�u\Q:_�R��*�䡳D� �Ɂ���L�$�W����0�˭e\��#,e�ޥĕ�l�5�\P��
8�Aб-oi}��9��Ϩf\�5;ţY��)^�8c�ȫ��o��A��<3n�����E\=���y��P�#O����_�5����I��71η�3�`�zlh���-�� ��G��-t���&>TM��*�|�x
��M�0jnL��m���pl<N]�,�|E���tZD[d�O���B}��:���'�n��t�'�U�P.� )ć��s��OZ�S�%C�# ݐ�v�*o �|���j%okA����g���< ����1�WO�\"/��s���p������1� @ҍ�&���CˑIQ�Wvb�V��}V����R��2�3�
$�t��k��=@x&
YNw5�Ű�4K�#���Hl
�^��Ϫ��مߓ�W�!Cx����dM�d�E�Q��Ⱦ2{C���8��͗�
�	�ΐ	mu!f#�.�:j�q����V������j��рw�j ǰj�ѩ��%d�T��^>��eoP�o$��'^���%{ʹ�͝�f�i̋nH��`u��6�����F<�l�!���#T*��7��ePjo��N[ߩ$Zu"�ct� ���+!%Md����u���=j���F/�rj�!���R��k+n=7�]��w���h�����B��G??>�5�qx�&(
��!.�	w��fyoL�j�z�Xʾ*�Z���n��ڝ������ෂ��m���ͥƦ��Q����x�mPu�[m��|\(>���B��S��d6�j��P���@�p��9�⽙8�>�	�������1��9��t�yGT�����LF��<7�i�i]PG��c�ݤ���- �K=�Rp�pK/Tw)HTw?/�QI�>�g�U��`�y8N�֬ׄ�[��ؤ��<�P�MӿzP^�~y������T�.~q]�*���K�'f]~�Je�v��#00KFоa�.y{zalG��!,��ک����G�����m����m��sh>4��#U-q��-�F����`�Ą����	�AꊒO=+ٲ¼ф7h'��i�nq^K�`�ܬ�K��e@�^ꑘ���ш�v���*H����,A'��P/*{�4t��*�;�hm�^�����HP6r�fwV������,�J�<.����}A%	�1b*��(���٬�c�B(B�f��S�P0c����l��7H�[��A'��'��	��E<t\C�Ѫ늭8�/��5	����2(�+�ڌ+_�
Q�<]smB�#v�	Si��>N|L�q�h_��	�9g�+�8��T��$����d1���O�\��� � ��8)s�0<�t�� �"g����*����8<y���Vn����_���̼f�>�LWO� D�ЍL���UbTҳ�d����%����Pb��N֕�`���pHk̠�53���f�bO�H���~^�B������q�3-�E�zp;���E���܄��Ͳ$ӭ��li�nq��<�����:�s�Y43������������=�����҅Q�֤���������65e��g������,9���%��#?�r��OF� \�������� �%-Խnp�q�Q�`����u�tK��6E��GOGG�V\����x�Q ���ҭ~&�2D�\��v����ﾢ�ǲu��9�Ph� �_Xt]Z�7�4k`Z��Y�r��{K��r4�
^����n�L���H�*#�� `lk*ᳺ���UV�ӄ��j�yH��������9�_�>/|�AǢHPo�-!�(��`�=�r��.L:.j��-`2
x��z�C��1"?c�Y��������LE� ������{��ٌa.���QŤ|�V\X�{Қ�H+1���Ay�#�q\����i��A56:9b���$o5l"��@X�V��fv%x`c��y��0��+C�}bG��G�x�5�-Cj�p�r�$1zrX��C�{܄��H�������8[���= .#׋��EqF�i���e*A�[�⑶���"5!����\ �4�E����X�C�]�o���M9c����ٟj�K�4�
����~���R�!J�ˬ��_<)*?̤1� �ĕ�0��J譁o�P]�6i+ g�-�R{��Ѻ�T�W���#f�g�cV��hE��q Y�BV�m�&HL�M(w��Tu�����R�]7㍱�����G(�"\���)N�?���n�Gb�sӼ|�����{2B�N���f���n�����F�W�_����cl	(�H-����@��p�
T�3���!����������s
�{�S��Pz��wHpo�\�@�>	?zZ�Aa�W���F[:r��S�w>�%	��/����l�4��XF�d�1}x�c�zݹ:���B/H�z$��ǷnO�qu��|�R���@n?T͕���5+"_/�-.����]�7[e~te�}�ww��EMw� ��Vza��nR�a��H���:v�A��0b���ø$cR�
%\�}�(z�O��\�ϱ&#C�CH�V��]+h�O�Gr���Aj�t�GêKմH]�5=Y�t���c�Pi䷼�|K!�����+�'��Jᙠ�P���=�ύ����v &���
	F_�H��r�Y�0�U�v1뭤��l�z�1�i�n�2��I��� -�50&��'ϭ�A�ߚȮ�rИY�Z���@�e�������l�R'lz�=��$]�a7�#�Cmd|kRFvB���Us+�8EF3���]��K`��@���ze}�VI=����d�#����%$�K4E��6=7`�͛A�f5�__�ޟ����^�К"Z�I\�Q"�G8�;3U�����s^����b*�Iͷ=�^=�5�ڧ�Zzӈ�܋o�Ԧ�]�6����hH2��Z�Ԛ�K��pI/� 
�E��`�Z���E�Z�]�WOʫX�ţ���*�*,G��`�B���K�&5�V}ߛ5���@얖�����ޯ�T�%����J�X?�|o "h�AQ��W�|���Z`��4H�6���J��п���x��Ѷ�lC1O��2���Bi��D��m��9v��0�y`� �'�UOI4k��_����땪�Q]`ͽ���[d�l���`�.f��3�s@�Hg���i�9��gl�����<R-�M��&vg��u��'�2f�H5�%sQh��BmX0T�[�\Ю1��&}}�\DC;c� 7�TUVs�������}؜7D���i[��jW��7���/��M2A�=S��h2/�	�&%�W�Vl2j&�n���\�D1�!A��K�I ���#��D��[�D^^��4CJ�
J�Px�f��Fn�76@���X ��=\��i�΢U��z|p�Z=�V���^��IsU<���wH&՚�ej�M��Ur7����-r3Œ$�n����MYD����C���A;.�[��vH��Z� r�B����IQ�� ~��=@���Ժ�Ya�F��f?6qZ�b��#�����K[�w�#{���C4�b�N*TѢr�����v��i�����]Q�9w�o���r��t�-BU���j�K�j���쑫/ c�?�%��<�1��lyw�o�|��/�/�qڈU�4]:27�wNXz�et�0�|�ssnɂw�Y�&|c��mMJS��h;��ļ-��%Y���8�Q���K�Qqz2�T ����|^;w%���C^��^	��3bTZU�_\gk��)CuF���Q��s�A�$++�!�v�#rY�A4�6QƧ'��;�py����w�PE�'��y2f�i�)����-�2Np���UQS�Ც�ޖR0_]H1�/eyl�'�U1�{���j��Ɖ��P:�����Fo}L���]��>����y����B���Wp��E�a��N�Zn?Ƽ�3|�np8��B��1kp$��k�:n��q�@e���Q�{��Dj�ﰆQ#��ӛȑ��䭴-����@$N�7y��Um"��э�ܭ��[0Q'��*�<w��0/�M`�����W��BX����U��R�j�bxj���'��hug*]���o*ۓ㖝	#	�^���: j����9cS���ۣHh^j� ��ф�nD&_������'�4�8 �$h���z��vg q*Hܖ�rJ���ud�f��^�V��KV�(&��I�G7�s4Cy	�}@��H��o�b�e7�QQC�L�����`�r=���T͘�ϻt���l{����j��<�rZ�WY��_��ϕ��=�L�6�E$�-�.r���Dn�T;7�SϞ�Q�*T��)�	*��W���W�˘�
Xg��E�2�1fk$��o��*F+�𪱺
X�Xt����gݗ��L�޻�13�a�qlW���0X8��_ɴ��?1_`�J�tt�ż��6$8�0`���ӿBzl��(���^�z/RS���?�W,��J_�P�}|ރ���Bǯ}�<���&�'2�����)ꐗF�m�D�}@�W�g_E8Xk�?/�/]D���D�
N9�ŧ?#C3�hɶ�����T]��$�7V.����M '<T��	z�
Z~)Q�k:l3i��l�?,̾��2URkٱ��a��!~����Ԡef� J��A��3��㗉8�6��b��W��*�ʺ���a��톅�]���I�7�$�`�Wۆv��Q}�4;�G�D�X-��\%Oxa��_
9Ah���f=��"3'n�?����[�I��K�38y܇��B��'dB8xh▾?2�?���H���(�y��4.�r��Z���%��ԓ�����h<2=�v��/�
;�/�ޭF��؋��#<j�4���y�%b�V�y61ԃt�M�.���A<��e�	�V�8��Ϋ�N���g<�$�����{�/�]3��&�A�?�!�
=Ϋ.;m���0���/r����SC��# �`ʹ�����E�?~@���o��� @	��w7pJD;m`Jp7��wC." ��{~
�����'�A/��Q�ٝ�I3�zI#zG�XTYvUj >���C��RZI��Γ��6��\�:��r�*Y!���Ҡ��!�D�*:1��y�EX�&�tsgI���G9���5��Q�el�Fl"��ᧀf��\��������j��������}S$���9g4����+C�lC`԰��*��S��G~��ϻ0e�ܝ�h�����,�|f��|,Ǻh�PN�Zh���IV�-g	�A��ѩ�t`���9�я��X'p��%��C]�n4��c�lH�_sM�'�R�d���b��Et�=w��LX�
�0�q-�G�C�v-є���K,��*#��1�1�����e�w�T�6{K�H3+�u�N:���Ν�2:@��m]n��Q:o	Ou�Ɵb�w�xR���?��p�r��F�~_*pm��ct��q�Q�y�~����۪q؝Cہ��h<{C]��ؘs�J���^�m�@����i.�y�6�&N��J�障Qm�s*tMD�<���P�H˔nj�e?�=H����P\ty^&�Z�&q;�
]W��7�Klc��'F�E�nq9J��J�&CRPM�O���p�aU8��ߤ�JsD������x��POp�����I��w�%g�poT"��TV�'�6�2�P	�YO��^lR�~AG���\�O)�v=Ts�:��t|w+��� �o���p��o_������^���hC�51�j'QTS���IE��A���<~����Wg`�����Uh�![�僧L&)u�r@������KĜ~@�^��/}w5W, y>��0��C��	�Ҽ|T�ܧM=P���l|���������KY.�7�S׉(0{iv���mC�@U��1+�į5[P��,�!�+�������>����w���=o�0K�V�m��F�4Uj"��_���ѕ{Kf^Q���F�,��>���F�&��������[oIҐ�0���.,�?y%�j���)(9��)`L4Q���臮ٙI��,$��.=�x:�N�����[2��En���y�˃H^}��ey�� ���7���sն1�'(�S���MIU��7w���%������Vqg��X��_r�A׈]O�� Ȼ��d��1`��<:��a*5H��ȝ���'"i��1^���R�j��U�gV��Ύ�f��,f���L!���e\b3��ě��X����a�`�D�8�^{E��+o���
 )v��rZA���v��2G���:6�K���0a�g�JN�]r[y������F|������{��v�`�]ܶo�iBhKJ�tEzuʟ�,ߜ4�F�V�8��JЋ�u��D���R|GQ���\S��?���N�'�S?y�ŧ�NT�F��9 &m���Z����2"	������0�o�c��������ﲻ�|	j���~��r2Vȡr�p.�W���}�����(�� �{T͚6�B�E�
 5uT'�b��0"F�u�k�b����hk�ɕ,���s�3~s��D,z�]�(�ۀ ��99��˘^�n�4F٪�0�.�"��wH�@�W�Ŏ������R~�#��-US�yx�o�wW�יx,<���e��0ÿI��v�!�l��rn�@����}!�렛��j=��RG��{�k¢�+ C�������<x1V�^�z�#f�Y��4tJD1F�"Q�*��8��	Q�i.�������;op���T��*m�\3�X��������ƈ*���LC�_R�L@%ф'&�sMl�0�HY4�-�m�2Z���Թ�p1���֜ѱ�馪��3?St��D�e���D´��u�
��je4�#�*����+()E3�v>;Ҽ�AV�����#(��#�ŀ䴧��Pb��Fq����O�ډ�����R�/IPvw>��_&i<O��D�HB���ۆi��o����Q�]��m�6gy!4�/�|����	ZJw! &+t�d(;�h������#tо��dR���~�;��/����c֝�z-�s'V^��&�Ey$FHJ�1���M�1���<bP7E��[(���k:�<���z�����u2�u�)<u[,�Qq;/.�;��+$�"w�[�,�
�շ���R!��������Q����X����Y,�R�`����G[���(L?@`e���5��*�Q�H2��޷�L=lER�J�krF��U�MZ�<������J����j�=L<*����o?G4��Y�
��9�z��S�{��������RS�!(SQ��eX�0�J�;*�'���a����/ݏg�� ��z�@ �X�B����n�0���E��
ݬ�=�Y)�!Ce�!E�q���8��ݏ�|$@�pA ۤ�QsaL҅�z�z�����RXL֥ �h���G+6�
o��=����!�m4��С��r����JH�����ZL)�����,����a��Į��/Xr���m���ĵ]Ģ)��v��e5�{��x�r!ש?�v1R���'���n��򛩹(�TT
|+,,o��_@�[�*��Z+G-Z?�h0Z����WQg�^^tg'����H`x�`|06N�[]�L�[�KWnA6,���� $��4/�̓k[cqL�5��e����'穯��؜o8rvu�K��KR�{�$IR�2��U��[)L�-9�-���
���iZuG��(����F�|���'a!eJ��j�;�.]��{%Y�f^|9�Uʧër�ǡ��JtT[fg��bPB��*:���i��`,�"'�k�mTڨ��2�8/l���O��у�T�(Ư�#y^At���o�;C���> X�}�㧟H��S��E/
�!>as���ù<L���:'h<���ӭQ�g��o��F�oq"�eq!�T��y7z�ޅ|��Y�$����M.�c��P�KkfT�{�\o.K� %�|_��a�Ic
�돳F�CU>6�����$��<�s�2 N����^��`2��P���S��f�m*Ol�+c{H���`�>��T�3�;���b�˷��vq�|N�l�Dd �B.�S'�<�*Ǧ��̸��ϲu�M��=+���j=�z��Ȓs���q����6�1�ab5���D`
f��D����^/U��w���� �xޝ�(�'A��q0������Zڪꍍ�((ゝ�'��-�������n���^ڙ��i<py"
S@���"�D�����{g��*>ai�6b11�G�@���9ĳz�P�(}���HPc̘f�w��]6b�(�1t7�˙�Iǉ�
^�8Ov$&�0~%I]JՏ��CT9��V;2}w�:+'�2��ű,:�x�2Yox�@f�,����o�9�;�@����D�<Γ�E��`C_�(�[�6�D�z�Q�������Y�J�����s����l[�ȵ�sԀ#^^'yd��]�ԧ�A'�c�˪��H�8�'/р z�i��W������9��" ����(�7�j������m�=�Z_v	D�T�N6<D�3R1�?[��kњDAs��Q�pO2�-���?h��������/w�R��Jh���³���ߊ�ܳr^|nԳ�� w��^�.��xFxDRX4�'|�Y	�p �	s=�hu:�e�k��w�7��b'é�S��)M�Fᕣ�֏���~>v'[�Ռ}�6I��z,gS�ga�R�n)p�Oj}%�O�Ue��'W�fb��9����|�e��Y�Ӟ'�<��Y7=�z��y�i�}po�Z3J�)�P���&��A��Q���Vbk�a#H�!iyh?����K\ߡ��A࿹.�U�9w1fC�I��w���^�o�Pw�+�2���n�N���ʷx�գ�L�M���ُ���0s(�B#|A/+�5n��q/��` R*�d��T���?~;KW/y��q���v������2�q�80ls���PԮEv��'��CN[S�N% �B�(+	�A��Njnr_R���to�=?!��9�45J�L� �H���eڧM��`��J�-V��`�=����#b"�E$5TЫ��Z�]¬��U��%+D6�K}HܴKi5<�I�e'�+�������Ꞗ���o�k��N\���w�fI��b�ٰ���L��݋p����a��ӽR�*G�j�bbFH~�l�Z#P{!1>�����J�Q�v��P!x���h<,
E���� ��t�~E�����n:�d�A;�C�oe:#_k4`;63����16���d���-�q� ��g��A�xI�C�j?����q��<W�{H�����E}��f*���Z��Ǵ&�0w����-���EH��)��'���n,A�(�悪�a,�/�0 )p6���z��ի=Ub����&pȢ�W��0S�0�+o��Ӎh�̿������a1,�o�p�4�M���"�#�J�Ӯ��q�k�I�C�������B�i^Ż���������M�s�LI�5���O�ݾJ��Ĉy-������3a��TB�'�~W{�&:q�J���TtՍi��4
���!���qU��w$J��޻;��-ǣ�q��m��d�8��<�R?Hk�%��.�9Q���c����K���yoR�]�C8��Ky� +jF;:C��mn�ZA����B�TX�]��e���d`7�%�!%y���-z��R��W�8%��E^ߗ��	u�zb-�ii#��R�K����3A�&s"�^0Y�L�Eֈ�w�(�X@�Y����0�[+`�`q�w
�x��b�~Dt�R�2q�9��6
�ҵ��o�h�n�E�z?G]D�	˲��wl有�����!�.Jx!XO�
��d��ױ��I[?��iQ��o%{ML��g�t�4�t5?�CE�mh$�pљ�f�	#���Ӄ��)dzm'j�这~`ͯ�-@�&vg�Z�Q_��t�N�WφEZl�p;H˿?���:�����<����V&(1Ӌ��!�o�v��)I�0���֡��]Ҭ`/S^��" ����_��ڜ
U�OyKh��?_��lF?aS�Z��U�]���5��K�*��`����Iæ���� }s�M��Ͷ�*�A�Tww�*;�Y� C�ץ�C�Ŵ���VE'v^����0?9h�?��1���������,�~ �U7�3mt"R�Z�`�u�O��7{���[Q��F��d��7��9�u�h%-�~;l1�fE !{�DZ�q���h��Y�v��x�3���8��>�����-R ������1��*)ޠ��(�����Y!�� ����g7JLɄ�r��0���#y5Ԙq���!a�պ��`G~��k�sؠ�2�!�c6�jL��i�[�;Wk|�'Y#�Q�n��Wr�.�O�O;-� �������|�����_�#��b��`r��nJ|��UmM�'6�;,�0��LaN���NAV�+PX��z98��U|�]��e���M��l(eG��R�]j�s�ǃ�#�;̺���Q��E�>J���#ζp���>x����<C,�n
�����aC?m����ٚ�:|�jȁr���b3����d@�7��sE��#��T�C_Cn���5�Y�]}b��%�S�Ƴ�� a���/F�S�<��W-Y�Cwq0㳢x���<[K�+�J�g���\\PM��)=�2a�2��0��_?X�2��rV�t3
�i2q�,�a��̻�"]��zt1��&�����:R(�{��Z�!�گs�-�6�y���������M�:�|����nlU��ٜp��#%��!��;�<�q���x���n��D��dE�w����f����U���6��#�ì{��Ge������)$����`�nK'���`3#KF�OJm�E;����/,FR�V	݄�\��<��X�u�?~ٓ���Ђ�uf���S9�����2��	����Y�Z��&f� ��W}�~�K`�8�ۅ�mQ|-�2ʎ8�O�Nqp-�� 1)��!�P+�<���Z�ҋD�������V�6h�'P&5��^��?�D��F̲��rN�:����}���
L��_�HQ�I_�s�)���S'ar�|��kPq�-����o����:$O��`Pp�-5z�%S��Zpat�Qel�������u���&���>�՛M��*B,�n�:r+�0B+�.VhK�v����Rp����~�����ؗL��R|_䫿� ���L�d?�[6�|���U��;_ߣ�pE���T�C&�[
�/:��&�0_@������|�49u��8I���P�O��KQ7�ͼmD⍙�!�\0U��c�r�,b�́��#C�"����ebJ<�P�6ߪ �#�A��^Z���vn��g�_��Iv9��n)0r��|�eYu�a��n�Xq���W�#�c����*���
 ����A��Y@u�@H �-/��e��jB��rd��?_���)���Qf��U��u���a4�j��{�Q�_ݕ���XO4�k�I��S�Ͼorx��.��e����&xsƍ#�#�<���W��_w�D������c�_7]QU8�򘜠@r9C��O��8!Z±�[ݦ1����8�5d̠Kƶ@�|��'ōer�\W���-���MP�lkM)8��z$�ڐirv8������$ ���s4�?��r��Ȋ��Ji-� ��� 3�I�}�B��h.O:�ude�@�_ o����0U�~��l)
�r.�(�\��)R�)��rY�xL�Te����Wv��$]�ﱶ�;!�jD2��N���_�r4��,^t=�T�t�\2=��AN_*N�pJ�a	�8��S�ߥ_=��KZl���;��5�ɿ�{t{	�T0�U�\��}
��|3��Є}��N!Vg��zo#;���ac��"{�r���>(�ЫS���FI�!�vf������F��_�Zܐ	.oJYخ�B�r.ә>Y��v�r�Bђ����2��������S��E����W`�X�7Kʑ�P(`O�����v�s���h�RJ	�h>?��k��Ţx�(%�筫X�K�eÊ����Qs/,�u����l\K�
���G��'�8�v9'�-eG���E�l<;�;_��oe4j�71�Z�5��;J����Y_a�{5�]�Oa�2iLk������ơ-�|Ӵ�5�����R��

�?�y�o�L�`2ƅ�9_΀m�ɔ��敭+�������*]��A���@��`�R��Ǩ�E"�Or؃-��o⇇���I�)��]&�(lԹ6�k��خ�iO�3�H�;�GABTB��۔�J������Q�,V7���0����n�tת�BR[�<7?[�@煮Xu�N\n��?�vw8h#�� �a��� ����I-J�iv=h̟���XQ"�+O����{o��1�.g������ -W ���P"R[�g��bɣ�!s����Y8�v�烏G�S��΁ja��!.v7����AdL8[K�B�<v
�Ζ�h(U�}2�:aG�#!a��m^c�t��=�-�4_��ȡ>�l�9cE���~_bN��L��mGe$��v;t?i� Ӵ�ِP�æNV��k)c�,����IQa2�_�g-ZN��?X����XY{���#�iLŤ��rx�=�YŀXZC�3y��K��w�m�1�A>�T'�����6(���Y�����"�P���n�O�̆|���H-���WE�m��N��N{�3}�o}��y��Ӟ�[׻�����=͵ �gҗ�~s�K�[� �P��f��ރ�l1x�y�u3Sr�a�^ЂC0��o��ęKL<�j(��ֲ_�Ŝ}��x�C&p��Bi*��%�}O��Rz�|�98��^"��cP֙%�{��2|�����ǡt�٪����H;��[Pp��V��D6�����h����pJ��o@j�����Ĺ�
}/%��n����s<�:!h�h'6ɉ�U���
�\���λm���D���UYI'���4�wfh�����cd�"u�j�Sŵ��jM�e���$�*��[ �R1�,��C��̘HxY��J�;GU (z�g�;�d~�Dl���ŨQ����S�4�PK�h����L��3-xmˌHe!������K�囙s�]��8�}v��o�F�{!ՎR4%�Vڰ*���� =a�a�0^l+�.a �0��f��:��$ȃC�A����yw�\$��)"�b�b
�(�I���3�7c��k5?YQ�q�߆��Y-.]�k?K(�	C_2�\0J�t	I�\h�����k/T��	e�A E�������9~8�,��㌜�^ky%8s�O����(�U���L�����m�ۇ�I��F�;;+���,=+mǟ�8��t}�J]�"V��j1]�hv=9���@��e�G���j?.}�����Ǣ0�.���항퓌˾>�^	$k���`�p��R�ฏ�$�m,�^g�?4�R7��lC�9�>i�$�0���p^��0�t4ж��b���P-�=�LZ���H>��9!��Ov�	���h�_�������)���Y���xgI��2aV<�~suo��>W�-=?RDIV�O�W��|������� �q��{C���	����I����Gr!ڸR�(���~U;q��1���B�Y�fw�J��h�B�x"z�����}+X�G�nV��$v:� 4,��ɴwJ\~��Z�><��;@��[疴�spzs�����Bʶ6�?�|_�x�+�c'3%wP:=᳦4���$_�+v�`��n���7yό�juG�H\��y����3p�����JI�6o��8�� "�#�'e:I���gE�5�^ϳt�h�pU�q{�#JrQ�h�h��X���/���3MG-�|��ǀ��Y{��m$�5�����9fu�Ĺ��F	��?�O���	�6�{��N9F�gE �i���h���"Y�/��{Y��2�۽j��H#w��p��U-X1w/��JR���EB�Wz�������%.�����|p-li�믮��r�@ieսz��R�y�p�J��&�T]����2?g4���3�L��=I��<8����
���:I:�~=Br����p�����
��̞w�"$\�͉[K��b��� %J,fiI�@�mA���i��\W�6�a@OK�
�#��]����akZ{z�+��I+���ko�(��� ��&�f>11��Y#w��m�(�9:������=�z�"��y;`�%;׺��Y[�?�ъZҿ�6�u����в��擊W��j?P�鲢TR�X�]�G�Ͻ�.s�rx_����=.�x�\�\f�	3�mC��`�n��[2�-1B(|��!fR���:�����%>��`i��UZY��QҦ�$�2<��rUn#�I|�r�͓M+I+g�v;��B�?Q}������D�m�ɮ]%MF�cdN!7�h4�]���:x%?�����5�l���~A��9�KE�h����G��M��"q���ޮ,[��*"�N���r��År̹���]� ��KN�������_�Ke���S�\�Gf�˺���b%���X�@��9���c%���G��O����H�3�Xٯ9�`A46*�JM���v[�]�gQ��P�`�@χ��8$��1Y��f��w�J��<� ކ���*�c�m�7%�t��#	�NRsL�x:D=ȧʝ��pm�bH�a��k���浅\����F��U���>�<�
��bX���J��Rr����!{s�w"��-�Y<�"�-2��{'�`<e�98����$��V%'��*]	ɖe���8m0��H���	��z���W<\��>���m�,�dO�PN��s�%)�Z
<�ѧ1�3B��H:���÷�_u`]�*cg��!�d���Gk	8E�Gף��tE{�:\G~���[�$T,b�j��&f����*���RD�8��)>�㳷�S0 BG��X����i�$#iQN�H���� �r� �3�U]�eP�b����l%-ʨ'�����C:��4è��-3DV�D@�g"<P"~����v(����{l��,��!���d*��u�h�5lhae�Y2c��]���P�l����̲�ј�07�80Y|�,IY;�Y�=�����e]B5h�l���%qvb#cw���֥!�t^���]�f�G��d$[�v��d2�+=�B^��������qDW]5D���T�H ~�Ƭ)�j�C֌�[�r�Vn#�0�$'֕�Էn+�9������غ�:�?�`󵝅ǲ�_n =*�d��� 	f����s�o����UO�p�ҿָ�۩ �$��\$���|� �KjBz���y[є(�`tG������ӛ�yb���&{���"�W���bO3E�G?����v3i�6�?+W��8�O�M�����Ü��yR��"�&��x ֥:�������K�n��hv5��y{v�X�
m�N�D�t�#��)^}�WU��rh��q�fC1�Y*�R��w6rai�Vk�?�o̒����V�%z�S��U�n��S��Z��C�α1��jj���xr`�$�E��5��B�&7p��&���C��O�K#�5iPl��G#)~�AK��o"��Ձ�-�Q��z���u���Ʉ_�4�+�؇����a��1���<�5Y�	t�K�z&l_�8\�80��'x��`��}���٘im�cG��u�3R��o�=ҁXQ�"�=�6����}3��+3͒�S͜�}i��=������Zq�]�Eg`���K/�(C�um��#ꌳy�/&�;-Z_�s`��z�p:�`�&����9Z�}[}Y�AK�T�	|�/�\�Z�f��ƄD���w&`(��m�q�i.u�Z�6����\���G)`汧oS���ۃ����w�������;����.����5���?~��<m��l.�M�^/Ж�qBj�D�ԔO���|� ��]�&�)��v@>r�D?���(A�AS���q��wm���zZ�R�d�[������j_H�Y&�}�\:b�)z�[� �D�Vc�	C,���>,C�ߠfW��Y����~i�ȭ�t[���w�r[�gD�12e#�}���7�\��.�2��MU�y��=
��A]�Z��QL��UW1���ӏÞ��%|3X0F����h�#Z%�H��<�7�_jq���#��C.3�|���%x�HW�/���vukg^��y�~���46�E8�;�Ր���üJ���`q�7,(P|��<��6Ԥ
��\��FcD��ț��h
'.{���Lӓ�@'�t�����Tа���%��'_��&��L�=(�7�g���FT{���lA�\f��K8
l�}�zY�>2�Z�c%��*���E9����ݗ,[.p �+B��:�7�]gW��kC3��Ė��>�ݳ�O*��@F�����o�&�� ��Q6���������ݕ%	�)@�қq�� ��}ɶf�"�↵�k������A^��?
�w�"�'����,�e$=:N ��G�`��B�x��!��b~��H��w��\{������n�KzsR2ʗ���tw�;y�?P�pو�^~2U�f���Φ~�(%����������Dtq�m�˝=��$�na����r�-1��A��.�ٚ�caiK��r�q���oO�F��f�*A�pa�%4|6G��'_�,Z��֬4��! Um.��Ҽ� m
!e��tMx�)�����^s�)�>f�i�� |�Rz"�f���*����r�S`���P�ԧ���c�ۻ딼2�[���ԋ�����(8�E��-2�CB�#h�T��&���I��d�y3#H�#AF���h*�����7\y<�k��ѭ:�$�7��Y��I�V�ؽ�!),��q�4�"[Z]F���]S���DB�gإT���k�s�Ne�44���+��j�)�B�_Nc؇�j+��~�vn����z	Kj�ԟM���-���_Cȏ-�Irf��:�ॖz,���{U�p� Z�ǔ��z�=&n�e;��K�o�"ak���!^s3U�����|�6����Vjڻ���?����{��|�5NI�7?G�Rl(:�p!7}�C��ڽ?*4�&�v6�cV�������$��ɭ�
��&�q�'N��W�
b��$�tgĘ�욗��)��b�����B7G�`*��I��9���<'}���v/�p%����o#`­�?k��j�nK��kX����K� T~XX��jS<�tb��ז+�u�E� ��j��:S�W��o��0�z<��(��P-g4S�M��0�%��6��V�>��z,�q?]��ʘ嶢w}}�p�g���#�3��y���ѫF���W,T&�A��8R��o�L�s�cT&Wj�G���6d���ml���f
���ɖ�,d�`�(#*D*�c좴o��}�fA㟲���pgx;��M�~+��!�f��1�X��0�q�j��s1q���<��4����f��	�D�j߰`�K�)�R+����b�G)!#��:��N���#��G���n���&�H�Vu\�� C�i�fTH&B�_�e���d��G���kH{% ��[w��з�Y��cV�_f6N���i0���8����5Ǆȹ��HM��؜��GsK0#���|��0�.��Бm���%���ۉ�� �o��Md?��I�M҆�ú��TZ-��f,�|�ΛS�e�9oB
_��(������4�S�����Io��Ov��=t:x�����, ]s��\���!�u�ᗕ��eh�p���G��p
Y�K���wR�h�?h�Y���W��@K\q�U��A�a�Ч|��a�VϾF��4��
K��gPI��a)ͻv�}vj
�H��O!��,����"hV"f�W�	c[�39j�	�Z��&\CI���
�	���G�gBfYU�X�{�m"Є��G
��T.-xdꎨ�Bߓm�|�|hTy!h& ��y�7/n��6C�^�R�@Y
�셩F�5�) v������`I�څ�B�ݓE����H�ǢmeE'���Mx�
���i� ��ՐJ��,ڮm���h����'7*���=Ey�IV�����|�R�%��p�1ni�BU��/��|iB����:sE��	�Rd��m˂�¤!=������ �T`�Y�,��gF�[N��W��/ː��;��ٵ�R։#��n�ϓ��\��ۇ�of 	4 ��݆�����rmF�Y�0�͋��������'漰"�C
����u��Y|IG(�
�ك�]$u���t{�W���i!Z ���?giq��ܳ�J��~H!��v�O�����4�م�>4k!]���RO�p-�%?�*���Q���D"�Ǻ����[�Y����b��~���u3f��1��Lmߪ<�R,W݁��#y��mT�GmC#�� �{u���.���7s*�6E/�ң oM�	x$M���$���C��JEt�^ׅѿ�:\��/k������?�+7��^��p�23t��7a>e��2)-�IHӢ�m����z*/���Z
��:��Z�6ë����������P2���T3�4�[B�n����P��76ZU��� `��srL; �7~��Z�[���ǭ|�������h/�U1�r9��6�@�{��~�ͯZ|֥r�`k
���i�}b̮�=���3d���e�d$ބ_�-��أ�A�o=A�ǚ�B#"JW�����a0�[վЙ*�}7�I�%?-=�~Kj^3�"�8s�8�kZ��;��-)B�=CH ������"A���/ASo�q��h�j -^�Q�-Į�>W���Cy_V^��h�d�l^.*��͢m��]\)߂�H����tb����T)�/[�8GM��Nk|�lO��&���p������]x�I1�A�2���V�X3��G�Ee���J���W0l�7��|�$gk0�	�E��x�f�Gy-5z��a�]Ģx����q���
@+�*����[꣺�k6� !O���vi�IZ���F���OǗl��n_�mV�=]ȱ�_�D���N�&/�83�1�������1ٜ��6L�����I��eA��ח�O�E���}��NV�HSS��)/�^����� �0r�U9-p��<?�~è������X����A��.'D�b=�� ��w�诃We�)/��inE��/��+Z!�7fKb|׌؍R&IU8�L��:�p�$�J�xT����y$�ˡ�G���8��;V~]MH��AU5b�&���T�.w�5�<W(�0LIXʖ.���w�y���Yc�Ԕ�N&4������L
���E��j��/>�U�$�t!��)�iI:������@�햲�C.��c/ު���q�.�|L�}�������9d�t�t鷯�t�s;�My;]�=T�<Vʏ(V��p��v��}[��C��*[ �J����v�����L�*aS�!���^�K+g��@�U��9p�!y�"y��� C�;����D�E|��<c�c�q����Z*��3��ͯ��5��G�0�GxN�pOD���k�~���=U��)-��G�/b�f��X՞��\���cЧ�=�=qe�;��ʏ�:�y"I�>�zv|`1r��Ÿ�t��QÀe�B��'1EjF|S�����k��(����U����e:M�fêu��7<�U�}>�grq2�R
��~�Z.�#���%&��=��]��𢵼MQw�p�w��L��{oM�7�шWAĿ�)��o�(2,rA�Ok������!�uvN'=�F���7��N�ۉȈK��6�Lm�>:@u65��^���"�W G��<n�6�5	�F�H7���˥kDQ!�������='�ֲV�׉�\��TS)H�kK#��Cv�(d�3Z�Q��\��;!���v����`���.$�"�����ȏ��*j���F��|Z���}I�Q��A�(.�%�`(A[pg�Zlp��j�hWw*0S��{JV�9��g�D�H_�����8�+����#����G��.��i�X�{��z��V���iy�m갆���
q[�ƶhQ����,���s�͈o�N��x���&��5�I��y���k����&H���'Һ}�A_"t�֠0�s}����Odk��LP�y4�z�0B����?k1Qs6�_��P�a��a ��wD�0w{�;%���P�kh���CB�1���Iu�AH�>��n�jk�*������lz8��;6�b���;�PW~M�t�����@�}�(�:_R�ʥO��=I� bO��x�@�䒃s��o�W�
��q~�[e{n;@�M߻�#ڐ9�2���M�;��EH��I?��ZIX]�	�I��|R�6��@���Ht���%����
`WW�p�
4�Ŕ��J`�n�>xw��0 "!#Z��7�aE�>���֎���lU?��(�������{~��=���2"%���}6�G�*D���e��bI=j3�����ڕMU1Lw�0^3e�����B2fL�-/��ϭDE�e����7�����/q5���t����q���a+B:�U�����̙c�LЕEP32	�.�Q�ɬ7&D9��\��	P5�=�}gi�f��� `<&�qj�}�S�2ԗ���I�^$x���h;1]	�\�"S��с�e�(���T9c��x)���R����['�%��ʀ軞�oZe2Z��>��ڻ�
7�t�����=
1J��i,̯ճe�����&"��Ϻ����m�ʿ�^I��G&-m<�#�/�ˉf������#�z��{��+,�H�Y=��B�sU���C�S�f�W��ߔ>���1�.��\�x�Qb{�4'h4�ծ���M�Sf��Ub��zy6_�K�&�7�.�>���V��M۬��thM�ܥ�qUa�Q��#�'.S =Γ)I�!<�Cw�3�/�2��p�0�����_�@G�HI����W쒘���@�%���I^d�3�rʴ�6_�9�Zc�L�T��>��'�'�Dqv�լ`������N�8�d#%{`l""�r�%��/����&��Ԣ!�����oK�Q�}^�5(�V��D{�G%��uiX���
�0R2ʊ�_��*Ae�r�q�1H���;��!�j���_�h� ���h�m޿���%�r٬�^p�
��)*�g�=�^E����"1D�nj2��=n�������L�\���M��K9rc�W�FmG�)~��zeQWw��1�����y�,��c-.�̵��"!������D����Ǻ1E��2��peʴ �Rs�����"ul�T&]┧�TӇr�t P���-P (a�)�@�W�fN�CQ���5�/o���[�bky�y�q�w�1�Jk3�X\��\��E5�$����,��/��A�NܛC_��}j��x0.�r�?7���N�TB��R	��)�UÀ��J��?}T�Ƶ�/F�<�D쩷�ܞ�".����]i*����++^�F���.�]h|�-��R~������}�o�a72�u*X,*^��2y/L���ʧ��;�K]1ش�8oXG_��-븽Es6�)�d~���{5�@���Ì�>�s��t��� �C�����i[�e�l�a9Ÿj�	�[�@B���/����ґ9�P���@}�� I�OG��+�/n�DTvq;?}̲��s�WiCCd�q]���*�	���W�����JMF�Tt�+�;�A=��+��P~`�����d�?y���U>���K>O�M^8W���-�ږ���P�ytmץ��J�5b�G�����m�Q��)=�vV��K���l�͓j��:�\.!�g�D�6U�'!���J��Vm��G�,<[Zw&S5��x��4����x����A�g���,J)��=~D2��yE�2Oy���;��c{�\����x)P��7�ò����wp�����6�)��R��I?w�4Y�2C",Y�淦��%�2��U,�Z��dFR�tF2Ą`���j��i`5r��6���3ܲ'OX�٣e���ϕ�/"'u;`K�2\�����#�r���'�ʝ��1�%b�od'�$��8h��?
��-�����������Z6*r(4�8���E3��S]�<��-��W��S��H[���UD��@$�[$`�̮X�y�p}+�ꕓv�H"�W�,,�����
�dh���8�5 �����r�����#BЀ����J�.L���e	�����_Sƛ˝G��D���K�1�W���,�(�fhH�Ќe`7S`͇	�"W��S�ɥ���,��'c�Hd�z��b�2���+N�t�W�+����]���FU��+�y�t���A!RW�~�*��spo�+a�bc]��� $A��Q+������>u�y<д"�����
�]@r;�nc{1QW���sPEN�^��u*u��J��*�vMLbN�O	���%BJ���Z��-ڨhD�do@��f�C�h| Y�J��-������j�=?w�����
�̗�b�rD;���Ӌ�̊���ń��0���+�/v#�ϞC7%|
_�*��J�R�񶦠X��	��"���p��e�y�㎮rcN���I��x|ſsx�=p������q�$r�Q>r����5��b*�^k���Z�B�x]����0�,�m<)�!�C�yQ��O�!(�g�د�a�vU��� n�S���/I���]��	��ؘx,�j�P�&��_o߫��^-m�w�#� R��K=��E��?9��:�1(BL�tG���H� �r�`��x�?|@Fv�׍��k4}:Ή�'������K�(��c)&���x���)��{��޻A�##-҂n`t�ʹ�Q��R���#9xM��K����%g	�M��Vt`��X��tn�A;�ӈD��x�
��Z��u���;#5����Z���0%ud�6a�<%�k�xtȇi+�Hp8�Q����X�ˋMwp'�PQ�0U���,T����98ܚ�+��S�c륺
��O=�A�k�%$U�_L:9����L���ov*�f:��]l����Vx@�^'�j���艆�VD�z-F^^<���%�yVݙ��Ѷ@�v>W -?0��~����iujX)a,�|�m��9��?>�	�z���ޛ� �M��)����\\�פ��yڷX��w�����3^r��PWuǸA��0o��L�I��d���fhKHb��o�Co]�!�7So��6>���%�L*����� ;}u$F��/'3$4���"\��u��l,t��!�PӶ���k�8u�)�CtW�W�6��j��5V�|H�~Ϥ��
`��?�H`b���m!���1�����I�\~���x�z_f3��4�">�k,/F��F�(�ќ3�(��+_E�^BE��ɅP��K�=%�8N��y�Kn��{\�ua����A1m���1}F�&���1)��� Z�<��,���p����^ny�~�a���)�=_�j�FM�O��@�<����Ϩs�5�5+�|w�nqѡ��2�t�#u��A�9J�5�a�p!_�d��z��o��2BOY�@�>2�-)`	�2�U�H�X%��q��ڤZ�|�?�;H�z���H���̮���>WMq\T>���S���Y�ۦLv j���uϻ�:�$ B����4�<�R\Wr�»��)H2��<{}_7qw�rE�I}O��4�k©�A�.-Z+z������s)�h�o�U����ɵ1�0��<��=�B�+���#��T?�I!�¼��,�;O���G������ٕP�ln�J�ġ;CG������[d������C?�~�媤P�H��]n�*5���^�IZu�h�<�n���%��^�މfH⃏����׊k�U�5�AcX]�X�z?��Rs��L�"U��@���z�܃�ʄ�^u{�J�P�n$����ӲY2�F_D�=����Y��W�X���6�Z~�W�M�<�z[ck�<0�	 ����k�;t���B[;��\�Vw� ���е�Ku�ʯ_l]{�Р@�����rJ�2D�+q��� ��b�&u�����=�2�1�ۣ�cFo@�}P�ъ���R^����OoF����t'�NJ��o�|��Њ��'�f`���7Xa&�"�㲄ܒ[,���.;�!6e�/�X � ��6O
kx�I`���?ݮ���_~z�I�[�H���S(:t��YpLMAh������Jo!���ۆ��8]�۱y�X���_��<?hY��v[�4,<��:���}|�| rd�uR3�wCm�E�h�`|[����,ǀꇀ����`R88)nh#����n��x�tO|�3C�eW\��p��K6+'��5�w%z���sIԺ�,�����@�Bt�:�&50䟈>+��H=�!������@�:|��<�rrգ�����c�nװ���7ɕ����t��;j���u���X��Iu�iR����Q�͔>0{��Tӱt��b���À�h�v��ϵ��$�Af�#u;�,s�����j���)�f&.�G,Z}\w���^�E�"p���i����m^��B9W�N���I�Z��M����#��C6�hi����<�{�����~�.LS#���D�|�����ȼ��X�l�Ey"N�{ �.�y>V�{�1��Pb��J�����q��wYKC�:K���</g �:o&�C+r�W�ڭ�ϏO��x�=�[G�l�z5����N�Y ��_��:p���3^u�26*�ߊ�UI&6��+u.�^�_:�*�����2t� wY�N�%a�V|	5�/�����ں��#vHSR31����E�~ v�g)���%sxy}�a4�@?a���Ch_hP�E�
<�"~����S��B��;���:b���՘��k8�_g�3��@F���ΜI�'e9��^�a1���)�����΍���_SZ���!�fg]&�)��%/O������|�b�3�[�?�*|P���G3[� R>�,r���c.�a�9��[�Ce��`R�K'�Qx�����~=���df1��62����(�!��:���5���� �I#��}i������O,�Bݵ�V2���&a'�]�0a�J�i}�bb�H#����<�f��\A�	;��e��&L�#������R/�>���?��4��㈱�m�L�GE+��J	9.�tl1V�FK�*�n�� �������N4P˘5� +��N^��CJ�v]�n�K ���]�{.���}��}��u|�L���������X�������� ^��{&��;F��Qܡq�τ�s������<3�oK��xN�]�	h�k����� )x�XB�S�(�; �S��O6�q�:t����eA��u/�rKL����7bH���;��p/�3GZ]o�$����#��Xh�2��4�'\��x�^n2�"���Ρ�8T#�z�!����#�E���r�#��Ji��,��Lj�+)Ԭ;\�:(Um��aP������S�EQ��6[��/��7���Yo�]�p>��ΙR57P��W�D����?��`�����D;�J�yu����Q6���a�+�fM?8�9��~�c�`�m�"�@�&��$c+e9�����s�!��,�jp�QR8����d��x��0!��ղA���d�T�y*�j��vB����7���t��U��qN�WY���	�����Cc�/�6�ڣ��c4���*�x�'�(��|Ԟ��B���(IkG�A2RZ#6ߊ��Z7�[5e���(���5^R	@G���m�j�����+}}F���+D���Q҇tI 5[
c�n�c.�jO힏Y籃������*XЀ�1�gU�G���7�J3?�ӱ{8܉p4D����ۮ&��|Uw�U�N��@6���g\W�R� Ƙ�%v�O��"k�Ͼ
�a�X~�/��';�Ux���i�ݴ��l�|��r�/���(���&�������S����c,���I�E5H�xF�-H̜{V��F��'z�D?K�E
I/?zm)J\J�ogtհ-E�<v"���P	g,L 9��A=q𺛰w�q��-�GZ��E�{L�A�ǌ���/��K����m�����u!7�s]���-���q=��+�x=�c)w��|��>m8g���q�EU"���hd���+-�v��4�lf�^~p��-6��(l��c�i�t��<��2���L��B~��*���kh /���A�҇��4�4c�-��<(�	��-�ޮ>΍�O��z�<��]'�|h��}�1��T�0�E�jn9�B}y0�	�5���h�ww��n9�e��d�r���FD��5`?o/�"���G��G�E w�{]��yӺ��d�ަ��@6��F��Ƥ6Åص��������ۗ�%��R��i��X����p���"i�Zۙ�r�4"�p�q�ZH���;<T�p
�n�S=g��(�n� B3e�qTX�К��Pt���[�O������ݹ�T'g![��E�h�M�Đ<�]_�7�q��$̠����VW�`	����J�S���/�� "�,2By#}p9��zɶ��
9��h�b�I�cۤ�:� �_�&s>�t����ȱ�q�=�F���>c�xh��5���h-,9�3�2�"^���m
��^a/��m��K* �8 �1m �S���+q�r���8�0]Hw0og�Mv���U��ҵ8y)�(���5�)^{��b�l4����lVx`e�]�T}��H�y��x�?O7����v�:�D�E���ч�J�_��Yo������pum����*���eM�So/��KҴ��q���p��e
����F�L1?,�<5���P��l�k���,����=��x1̡��ט��x�kSnEن��h���!rWM�����������",t��'�_�K��v5�	��q�a�|����m���X�B��2������DN�C��cx�/���2��
����O�S���[(�Ɲ�l���`�ccLh�@?�ٙ� �%�$YwͿV]�̧kR�	���<A��z[Xm��������'!OA����P�8�M�8�b���{H�#A�[op�r6T~�Ȱ������3��	��?�Vm�����p��^��q[����ˠ��ei��[�=��a F���:�b��`������0s������A��ײ��Ë��=W�H����/q�ݐ��E�>^J�+\���%a�ba���9R�J�ե)�Sp��yPMv#5�}*.������Pe�@�����!%�L���35D�!��&�D���)�~�!�^��W�p=�S���#��l�H8E��Lq�fi�D]�(�Ci?^�n5��"o�GYW8@x����x�=��ֱ8�6Mjvss���YG}��k�}ͼ���\�T� I�gLnf�c�i*���B��SPǍ_-P��hwp��6�$춽�4�Ryk�#�]��q�� �oO��B��R��@��1BT���ѧ��	jk����~���y�Ҽ�):-zkc_��B�=P�؊#K`cn�Y�?�[��uV�g�i$	�|"V4��x�#D�t~�B�(��t ʅD�y�֎�}��K��'�5�9��\�dGҎ[<m��L��'/����md�F�2���:y�A-N���{�MaO��i�	���q7�t<Nψ��z����{4f�C`x#	b (�����	�{��0�m�rX<_������K��C=��H��d��l���R6$p�˝�bRh��l@#h��d8�/�rs�	J�M����X��X� ��;��w)����/�)�(a��c@��1�X'�����Y��0��xPLۇ�� &G"8��N\�uIr�~������O��k�(�il4N����+�y��?%:�������r�GvOA��f�ݫ�j}��<R��B~Q\����W�ߥ��E'#Ao{�l?���k�	��{��.H�.i��z��ٶ�ߨz ��a�"���o%ǔ,IaIT�>�p�d�#gu��7�ހ喵�0�/�5S��O.��؏�����&�����,��J�9M��j��j��tY��K��ڑ��@=���'�)�ư+]�7�E<D�����+Y����㔠E�U���W'+3���ruȸ!��b�C�k�M��)��6�߹]�S�����)k+[�*�"���'.�t	s�w�(%�)l��q���Pɶs�_��-4G�֟Y���;|Aq:?ž�8��װ����vDTة�R,��$��Z�i�R�zu�ܟ�a(�q!&T�Kf멢op:#�-��.':���\����������7Ծ5�g����MITXI�W]{|�:�7�e܊��?�[�=x�wLj�LA��ȉ���
��7���)�0)�!z�YH���7���S>3�&� ����n�,�[j}�$�X��j��
�5?Bp�~��T����5g�f=^��cj �4�)P��N�w��-��傇�}%%w����Ŋ�#�%��[-��:�	>{�5�b�����,��B�lT��8��:&��i��n�D�܈+LL�|�B����fgc3o:��V��R�t�;�3��_��V==U�11�a��6�
F�4"y}�Qz���%|�x�\����*�3�û	���ǔ���W92���oS7�pRQ������&~���P�1 ����H872�4Z���/�湙�4�M[j��Π:ވ������=������j�[%��>+KA��m��`s���*�I���`��z�y�)�lz��0�P��O4�;>���`�MơZaN�Ȝ{q́��n���ٝ�����IXO�+�>%S����v�����z���ĉg��ߡB��b��ߛ�ٻ{����}?�N?�S�d��k,7#+$�"zû�b�]Bu=�I�|�N�"��2��A�������;w�32���8]Ѷ�
=�8\A !��[�3#ĝ/Ӧ���P9�c�r�p��?I��d�Og,[��K��$7�e��� Y�T��S�w�*�[���z3��ld���G����Adx��lU4����Ёo��@a�y��vH����A�r����i��yz���TVHM���M��$ ��[h1�?���j=d��$~�	�pr�<*G����p�*��n����8���q)X�ø�_��:���sPŀ��(�������o�wܢ���JC���f�:�u���^�ȝ�|�S���X�yɪ����A�rr�C$KMGXҴQ�� ʃJU��������:�F�;��U�ͩ�H[�P��U���2+jʖ��6�q���C�*k���\ma�q���%u�d@w(�T����L���R����?�@7�'Zl��"���T���i����b���K�eQ��{����ၿ-���^�@�� �G���i����c1��F��AW�g��֢ٷ���D��e咤^���А�*������,��;V�	}�
@�� L�<;|;��R�X�/�?ͼ���!d�+�wA�)�q��v{{%E)3�F��q�� �/���τ~�~����2Ep���c�q.C9�N�NG�5�cV��8�w@-�?�3k�A�Q��T�NiR%���aL��	�ь��; �-��LC��v�����ah�4u�<,�jH�[�h׾�A	I�<�������]��M�6�X
�O����]��}��b`㫣,v��E���ŷ%\��SV2V@F�ׇ��[v��+"�S�Q���pS�qu�؊���6��Q��\�N\�Q1쥋�]�D#v\���`��C���Tm6�m�X��ҭp����'������������1eV�ѳ��X����"$+(j}��I\&�%�����-��JܗS��ʹ��3|IPV�l��BFa��6R��3>�\�<n������菷M���2J�M����9�7F�������L��m�T�����StZ���E���>������QƨzZ5��W&8r<����'J��	M�KxMD���*���Ao������e��/���X0ӽ,��ƛ@�	X��G��K\=b�{�
|���E��W�΢-q��ֿ��9�yц�Ш�uzi���w���9�4J}&3����Gi#�{����4B�#R	��],iF8��N����i��;���CƂ\X0��pm�'�Hή�p���͟:������L�Mk@��<_���49M'�e�s�#��t� ��g
�f�q�oZ�^��'���F�~y} ��Ŷ�6t2)G@q}��b~�dˋ�
8�S�?��8�}-#gΡ)�$��g3B��TP��e�[���G����GI����y�*Ɩ��ܲ]�]�{����Y�x1��r����8j����tb�f�l��]=UWxy������F��J-��|߮D�l�&� ��#�'��?!EF�}�?�'��������VM�tZMX��ã���V2m�6�~|�O�M�$5G�jt�R���a��r���_��?=�=���"  �p�����B+��c�\ě�u��|2�Q�g�4����^�6��>��R�ه7Sh9N��Y��C�c�k:��ȓ�$Jj˩��u%Q�)��e�g/�[����Y���u���,����VxT�f["Ti�D,�,Rm��(�j�Xǥ�+p��(�,Ө^�6�V �� ��� �w/���E����FG�2�J�;���Ǖh�#���9N�`�~�t����1�V�&zp(2�˞�r��A"D�d�^Fw]H�M_
���${�4��?��#�}���[��G?�RYM�J��ky�u �y��vh}���`���1�^n9Q��uB�.DV��G�ra�豗����
&�G�C���a1��է�����6{Z�\i��{�C��¬�	����n�dEV��J7j��^��E�)$�حS ,�n�+^%�0Y&����)� ��\#] J�˻��yS�����%;�;@͓;���Ԓy6���kֺ�Ԑɝ���@DD�I��y��9.�c �3F�a�� K4��;��ĳ�kcx7IG��;���mtʥ���Y-ƚ8p��h���ޓ�j��g�����nٹ������0�,NG���_ʁ�ېI��OZ���B������W���	v+�s��0���dNg9���P�俌��_\T�ե^e��l�h�wp�{�p?��B�#�p��].������J���Z?ǀ�q�E�M
�l�>9�!�b"�����s��hB)\�|3�Sgۯ�Q�SRv���I�G�M�IT�+6�;�И7w��K-:`���)[l�|�G�N&Dr��?H�X�9*vn���܊%�Q�o��Q�*F�ۿҀy찇��������#�͛�{��Gg���+1�it�$?*�O��pHp{�z��X4n	�
�N�z�P����.���@Y�]�x�P�����3�;���;��9t�0GJTqǤU��m���|H��R;��L�I������h�ۅ�of��ɦ�+�n�q�q�
AM�)DP:i�Z��2����ܳ��EP@�v��S�J6�����ny�o0M���8M��ne�q��<�rm	�<���t�8{q^�D�yJu�<�8Jd�O�]�b^�m=P��h�ڊ{`�eq�+D`V���+�v܎<s�2��3��)�~��.g����{�Y�xG'1����,^ `I�Mp�U��-tݭ@]$��G�/��M��Z�3 �&������)z�x6�;�?n�-�r��
������.*��]�PP�1�ŋ�s��l�|���8O�Z�m��>&�f1 �pQh+��ʤ��9��U��h
�އӓ��'Ѫ�Q��˗�(�I=��G(��L�21"���nfC�^����Xd�êG
�T�ْGz�
�K�=�S�5x��I<Lk�):]rz��[�!K-�<���sr�F����@��Ō}D�c���V��F��mn��`��x*����;�=�3E��b�����Ԋ�Ձ�v2&j9ck�Ll���.��
�-�:��.���iL`�m�7��Aj��1{W�����*��8a1)h(�!!����=����O�;1vd_�k�� ɒ;��1��	Nw���GyS����w{�uB�s��?Ӥ1�7s���YB]W�5k�t�rb}>9�wlX�W�&�<� �z^GK̨r�Y�$�:Q
?m	5f/?�(��u�W�Ò~��,�GB�y'Fz�%r�ƘZGR�~�S@>�đu�?�.+��n���zX����˥��'6&�����O����j@��{�@X����<�6�7�>��B�<�?��Kg�>���Ί@���!ݍ���� ��̛����`��3j��:�ʤ�K��Gwǂ���6�i�:�eo̵p9��,��G��Q�B��Q�bx������$1B��鎲�4D��B�	Rbq<���d:`.��x�<n�;E�L�q�ij\�Q��x���&�m��Yi8\�Lڞ��BҦ",�0�������(���5XX����Ht��k�{�&$���8��G�%�O㻙��,0"���'z�>��Kj&��Y��w�����Z@><5\~�-7��o/�?�� "Z�W[�5;��BB���F�����٬mb����]�-�xv��Z:7���uy��a$�D#]�ye��$�_�sT{n�	͐�RӦ.�&����K/1k�)�n�u_�N?!��l��5�)�M_^qg�\��}�`^C�Ƨ��<���]���I����bQg���}��7����ƌ�H#|�����@I��mMw1Wrز�L���eG���t-�t~�[��ps�ߘЪLI���z���R�57��搦&P����!޵�~�DWT�ۮ�[9�>��`Nt���a�
��c��N������+���*5�+-~.��l�(��&Rk,���x�o>���Z��H	u����H�C�c�EU�e\E�䛖�b�ͦ��KNXLL~�nX��Id���駵5�ri9��m<R�3C�lް��
��1�k���dI�K�!:b V j�����ӻJۨg�Z�8��e�}\͝���L"#�#'%c�ך��sw̄<�eI���l��i��!�Ke�!�5�O��V-9�����vܸ�ୖ_H�U T��i�_��ӃheN�����7:@rm��������T����	�	��XI�x��~��q��b�����n��Yq�6
�,�ܸA]�T��f��_H-AՂq�nv�9.��a� �?�E]�9w�r~	�;6V��\�j��0�s`���6�_�*���!4��jO#l�͡\�?��(�Q0�cd-�#.���n��t��PC���ݥ5N8R܍@vO'D3��X=ea�A�DC��q� ;��4�ǖ�p��n�NE��[�Y��=?��/e��.�>HN��9OE�Y��dˁ��C�#T74�W�v�2�u66nHG3IH���hƓWQ�<!��Bjn�wf���k����%�.���{hgd����|��uA���
�s|��w.=�ΪD���-�+O���B����e�Q�f�vP���̻����3\�����V� LcU)˭}f���u�˞��f����^�̈�>i'h!.=^��g�T���G���V{KY��"jfZ�|�ꕡP	��>�Vڛ�/��n�vɛbh:i�EpG��_�w^�O��(�߼�!��T��Fh�.�Us�|&�0]F��fl�# 9m��V}�5O�'��4X�y�6#��a��$��h%��+�Ⲉ�!�4�Z։`�5=�*xvB�|�2���@Ε��g�Y:�Y�L��bᚘ�)�uAVÂ���?�q�Uv�&E��A�ޚ�R�P�?u�qe��"�p4��%�����|���L���)FQ��4���Qv���M潖��o9�����"��S�� �'5��C�>�>�����m�}��J9G���X��܆��t��X1�$6�L��a��R�(�6����|A|���֙���הK���4C0�?k�I2��#��RY12��a���En�"ne���j������.Y�c���KQ�\�2�T&��ڬ�i���P{�����ݗQH��le����h��hԍ���%�$e����	������1dh���=�j>�ܷn�F��xlу��%^}��3!iI"��g���j��VG������2A&1��3c��W���yRE�)��|�H����Lq�cm敂��*�-,M,�B	S3��l�@�����()H�Z�椠W���.�3�"<�Nd��p�!�`g+%��f�D$�Qf��/p��'r�FU	��@b����No[G1��鿰ȹZz���Пp�o �9�;��F���G��$�f?K�-���9�L�O���l��߂d��DP�Ȳh2���?�}�h�v�Åbɐd,J��Z�s���Y��Þ�rf����k�e楩*�:�8�op�mL��4���$�>{�$
��8��'��j��5F� A���O��8-튱6�����w��k[E�EV��,�0],�����'�J�g`.�(BR�L���i\ ����p����I���_1�f���6��8W@ڽ��7�и�w�ZK�����Ś^4�:lo�&M�X�-�����3P��0�,#���_m������OC�)OZWۆ��l���$M��;~`)�Ҩ����	�yx��fz��浉>�D�H��
��dP@W��6�]����F� d����E[�5��۶6���ۣ�C���&ђ�W��������&��i�a���DG�`j�~�I8e:H��u�Yٍh|0)O؂"A�1
xYp�N�'���tZ����TN�g�	x����٤�N����0&��s�Hmw9�q�r+���ΧeR�z{X�B[ͼ�{�!Ds̙��0.+Z�(�t@�T���2D%��@�_��楬�c���;X�2�ɶ�����D�|���3�_,8�����MT�_�	)m�#����\F���YA�^6���P�d��K��4\�/#\��
O0|%[��m�
|T82�ָ�Z�.��6hX_��GPVbP-$��r:���O��~^?�q1m]�!���v�Ȣ 5�����d)+؁��$�� 2ł�E���)�5N7���K\�f�QCQ�IKi�T0�!_�_�[�9I]Z���f<��7"�;`������Eb�D�|Աö�'���W��	�-9j�#	�y��L3[$"�出�1.X��iU��ވ�
��r����<}��/S�b�{���9z̤g���6?�+�lNJ(��<�F?���I�~��#��`!��2�Y4�BZ϶߁�>��?y�Xmr*���_�Ax�o�Pbd�W�S��.���P��2�\P�ߎ��^*
2�s�N��2�g�4
U�THf�Sm�r8a��0��L�d�M4�>����~h��&������d�2bݑӻ��Ji��R���:�PQGbX".L}$�a���cx�Y&ڱ����rby�~Y$@>-�THWH����f^������s !{ h%W�K�p��Q�>������HIv�~�� i���
f���"�`:�麰��I����>p�\�J#?j
�?����=��~�=����/�ВB].9I�T�;�����E ��sB'<��F�ӳ���̍9��2g���nZ�n.p�rPvQƇ�t����%uZ��N@9�w�b\4�	��/�TU�"2j�㣕_Ɣ�^'I�)K����������1%'��SS�J�e2F术d���r^.ϠI�7_ȵK���RVX���SH���ƚ��w2������	  |��4��4�d�l
�`�.�"� ���zV��=<�&�V��c��O*J7ǆ���Czž��T "�])#���eL�TN���sCN3��I:�@�f���"\�#���]���'���?�5��k�	l���d �L`88A ����{k ~e���s�9�M#���7��y&���&jB.�rz��XCUH83�F�TC�m�8���l&���A����"i��=��x
맼�t��w�fI��M�26aP8�NP ؟��6^��?1����l�����ŧ��4��s�w��Wcq�qՋW�".6ê�"V�	>P�¬�P���Q�>�<��hi"T*���x�M[NU�w��-�<#I׽�~Z��2�`QE� |ε�;S��>U�&�Bg �&L��?���2���hO��s���7+3���&�	����EU��׶����FS���'/�:�[�O8�m�+Ӕ�_7�x �e�5�Җ=�#��Nz]��f���0��[ޫ��g$2:�b>`lP	ͷ��C8�,��Irզ���~&�ē�m�e��_�ü��VX�^���?;��;�g����t�/�5�����/���Q�Pc[Q4���5��%�x��"��F�{�
Z�=):�'t!ĥp���3:�� 5�a�1���SdР�V��p�i��(ҭAۚ��ª�O}�͒������0�?��22�N��>m%%_�
`���:*���@��V��LM����<�U��J��q��2��f�\�v�F�d/���ju9�G�~܇�^g��B�%����yA�
��7X�l��XSA�D��ĩL	}B�e�q�U����\|�VM��#s�lb�ܠ,���Em�׻C~K�2u6%��xu�]��~�l�>��Zn'�k�'=J���MH���
Y�������T�"-@�Ǐ]pDe-ӥ�H�G���P�����>e�d ����E��q8�0]�C����	W�v(�+��`�*����[�3-�繂�0���%Zz��Ho�Wl�S[o\���d�;�=��Be����H�!�O��UWh�!q�s�M[P ָĚ�S��I=Э�
�ё���8,���^g�h[%�}͉�۔;����X�(;O���vyzb��>�����Lx�7�l�\D��
�3,uK�a��\���z*���(5[��E���f� �B� #D��Nb�c�,��]���~Vm�:#p1v������C�A�, �\雤x��D�K!�r�L���qi~�v��=�R(��{1�@�G��#�j�̓�	^�ƙ���9�?f4w�з���Mk��M�?;n妷�zO�l���/�x�q�������e��K��/�
�R��aw�����.� � y
���&����ʗP/���/ŦG���"F��!"�U\�s����ȝ�����X�=!1w �]NY˺p���:���4�%��+g��n�~�ߞc}�Upv �9e���������Q�&~&��{"k�Z�jW+w��� %U�ع?���~/����� ��_��J
�ژ�L���|�lqL�cC�{��]\*^�b<���\��	dX�㵃�A�ˤ�A,����a�VrA��).!)�=g��R
�wf?ׄ�U�� TQ7�����X���Y�$U�����9P`ױ6Q79����em���&�CYcloO�W}u�wao+�V�I55h*��g�u������Nd1��`��5�\��c�/y���1 �M7�ڋ� J�1�m�*Jǌ��
�<��8-�b��⩒(ʹ[�\xZ|gbӾ�O����	�V�b>�2��Q�l���:�E�$#�y>��iGw��{N5��E�%�H����t��*(~�w����&��<����T�3��<@(	z�t�T^�T�����Sd{]oJ~X����#j Tyf�i-4�:+��� �ɩ�x=�E8����K	sB~�r���T[:�|@��[ƫ��Fl2��wp[!��q�U�����Q���o`,���76{im|QY�<��$�y���(��-����|����d���[i&�5.�5<���ʾ�+�@�W��4Y6�jؕ�c���f�FX��M#�ֹQ�mmӊv�c�X�VBT��`��:u�w%�4�D�P�w�(Tb�}}t���˻
��zO,���&��Ey��8{���"��TE�;�?j��o;�C�w4�>���2�P�!�T�F��I���A��x�:ߒ�yԳ���n�
)�eoHB���2aUZt��R��"\0� �`ȫ��L��X���d�!�o� �yi�9[W�@c��H�}��m��hi�y>����o��1)�M���呚F��7�����4>Y��.��r�}r�jfcd���0��(ڙ$J�s�ą��W	#�'Zx�����)�QS���p��_�I4:��4��)�L���pԝk�w�<��?��{��B���?�������#;��F߬۱cU��ͮ��S���A�V�W׷��٪��!��������K.`0��"��g�j�o�8{ө�}�����1��<P��t!�&6`ŕ6���|��Z�#��,���׎!�_©�S�|�
xႜ�n�B�a�,�1���S)�w�(r��lU�C��h:}3-)J����)FB�y�A�S���_����a8�ȗ�-�1ϔN�4<�<��0u���~�z��� 4u~ߩ���]g�Z҄�_ys�|�R�"[I�t
e�Hm�B�A���J��M$�/�+#����] ?���btd�v�{�}cU��?I/�cJ�NHF$Q���_M��қ:U
�(m��v
����n�T0@��Y�%�0��� ���Եd���և�cr��x�� o���"�bﵽ*ɇ �e�P!m��+�f\��_&�+	W���m�����Z�����С��L����};|C��k�ErkJtӓV���� ΩN���շ� �Z��5������M<��UO����k�sغD+y��Mk�R��Є��T�2���'�^��Q��_�3F�u9畛Ͱ������꨸�껁�L�.A�Ɏ:�".NaH����?��4�n]�3_̎"�k��� ��$!om�;��ZM�,qGe*U&��"G��%cUhG4����ikQmٓ\�@�A���uT,)�<=�G0q�Ƨl��(�1���ٲP�ߋ�W���RE���7:�?Z儘��eA��_!v�}-�@���y@�d7X��͜b�����Nں�Q7�\�cN]��DS��$�P� q��\m����v�ЙƜ��.�H��1V������C��@�!�;�i�ʃ�rm+)oG�j��"�J(�0m20듀���ep�-_��%�U�Tp�;�;𰌋����*�u�� �J��������)�t��ǰ�%L��6Ě$o�lK��&+���AʾF�0���Aս� �����ueU�f��n�b���=:�2?��J�b؏O��W�+-\;+$��ʜ�.I�.�����q�v]��Ξ��q�M}���+ၤ�C����ǐ�+��&6�V���@�����Àɝ���<��^6�&�Ћ����1\��b����<��t���J$�:��Oe���dA�O�)R�=����-+�O��*���qN�]� ���>B��<�^��y��jf'}NS��	�~	þ,���"&��E��@Aˀ���#?�[�LR��x�#�;�#H57�B�Q7SU��2���p�e�k�W��hu�iM� B�mO������.��c��Z��yᅸ)��<��=�7Z���i)��MnkY	�R.���0�ى�|=EZ�1����;5�gQ]���F��!��6\�3����'��	��+U����1�tD�Q�}�a�0+���k}���Q$�֚N/\<v�)����b��t*~m���:�R�K`��v�l�U��-���E"��z�udi�]�lp�B��rD���Zo{8S=�XOM���xVc�`.k�Rg=�q�H���#"�%����^_���|6޽�J�ڟB�h��Y)+�(�&xH��VË�gyP�;[�
09!5�09��b(���'g�t��HV>~t^@�����%.6rm5��1������1��Q��!��|�
hc�:�Qq��i�M�Q��mi�+�Ó����{jR;8J:��ҋ��T��3�L���"gHg��*��db]vO��-$n�0E���ۮ
{��2-$����V�T�R�hX��)����[�����\Jߕ̀�i{�:�G�*�3Y�&�?#I�
����$���7���*�ʕRh��P�0rq��|���-�.y�$�¶�,1���H��O�"�o���$��d s+.	T���y)�玽[��eO��Ͷ/�����P�tȘyU(�o�73�oVQq)�ű�g����4ۍ:�=��������|�Dd����c�m�cy��_є�׾�pL�L�J�ې�?�3d�_J��#�x�D��AM�J�����L���Oa+	�p�Bk!����՜o��3!�Yan^��c��F01c��@p���V@)����
$� �����dn���K~G�|yO~���OO�����n��N+�g�C�
��h��VD'q�@�U���f7�D����"��jԇ�P�>���^�YXx|v#;�h[��pL����1ԯԑZ�q�%���0Θ90dg�T��-�o{AQ��sFy���6_�u�va�mh�7{�`CTc�r�.��ٱ�����M��%���0��^�6�E�j9���4�Ӧ��'4�)u��Ec�h}m-�=����T�,�n���=S4$'"�+=H9 ���gK�`K��^���(
%Z��<�O@M^�F�Gq��p]*>�D�S8�`
z��aO�Yt��<X��B�s��/n��8>�w=���
���/=��ꁎ�-X^�/���?/�@C�n��gW�+�e��t�h���� �S`�? �ΊH!H���<��{���PZpſ{5�����E�Y�1Kt��;��S��,��4m��ZHA��v���C�
�E��{b��Τ�~F��mҳE[k"�j���<=Ƶ*�5�;e̝�E���:�[Q"4y�?�ũ�q����ۗ�ዢ_������J�G�;]����9˰����g�M"Z�
��np'�5��l9s�0	��pڑ��a�j@���7e)~TF�p����`��V ���<�t~"�ܓf�Dv��$���-S��6usD�ت�	IYk2�q떉�{-�y�"��J�6Uv�
���YAy�u�����Ը`�w���Ľ@v}a��a�
���=�~,CZ�
DL}kj#�&�u��F��#j�Au[9�֝�0(Y$�x�z��KY��qi����ط�m*�,��+��5@�/��s�ʖd�8Bէ^���؁��f��a�P�_Տ�#�)�7�Y����z�-��f������C�X2����06g������vq�s���iRʙ%,*�<��x��Q��I�6c����`;aa���6ld���O����SBL5�>�0��>.T�,�¢:��	���9D��h���'����}�?�m49��Bu$� ���� ��$��Zz����)��ђLuM�	j,U�lw�-nWl���`>��\i>�WՏA�a�P���ۨN�����3ՐB���o�"Z��A�?e��;��)e�R��~����b���D��/ {iŽ��􃴳���.)� ��w���	���p�E����)qKoOs�;�py�尞_�Щە��G����p���*Qy~����}���n�i��?#�����]�7_�A��nx�4c1��P'T�*�l�o����)-��qZ� �+��2ް�����*�]Ģ!�rj�u�hNR+��u�/��sɍS�e�(�Vr7�:��p���@��,p��4���U�<LO�]U�<��e�H������Y�T6 ���k;��&�m�L�S(��7�ǃ7���Ly��S*G����,�G��!l��������o��Ƭ<��g�y���oг�d ��i�r7��v��*��]|N؀=M��F	���l�8�:�xks1���h����F�%4�r2�k���X����^6���p:�@bЮޓ��\�8H.�T�Kb$Z�[��o5���|�|��*�p	�䌡���t��j_%F���VRn-m�4Q��J�-2�N�.X����=�YL���U6�U�k�/�
H��ߧf���D[7���z��Q�K�r�&��U `#`,� �<-�$"�羣x��P��=��-�q��RQ�8{bo��ӎpЭ=\��GE.ˁ����!}�'���*{��+2�E���,:��Y�;X�QCZ�&����x���"�9��r.B��$ D�����[�Cď�d�(����80�*��{<�c�A`�U��y��y�ngg3d-T�����af��~��Ω���I���vN�.T�Uj����hu���#Dn�V"�_`�	1�
����&�9/:�����Q��e�c
���Pq�x[�s�Np`J �Mq�Z	Y��Xa��d����WS.����R�qyݪIQ<���9�~^c�LSN�T�������+�aFp�
�����U&������~bR�/c�sS�^�wV��_@�E�a����
�Y	�|{T���I� �HC$�w��DN�X	)��+�w�=�AХ����ŝ���c�)��)]�I�LӐJ��.t��Mν�]Le������,Wk��ġXxw9���&K_K����1�+w,v��v���G����@+y��t8]8�S��yZ"�y�g�����y����jL_���K��)�����26߄���W.��1M��t� ��(-k.g�P�:�5��?�y�`t9_�h�M��El����Lӂ���`d���¸��-A|� x�@~�+'��!�����o_�����GZ��{n8=7��:�G�yD��]��l��Xa��W��p�w,=�R�]yki�I�తo�%`7��ߡoQ� ��Q�)��3�R���
���n�A>�-�a�����=tOQ�'�/�WD7������+:,�9
]+^' ����񍳡����b'Wַ=D�7CxU��.6���g�av��U�Uo�uΛ��?�ڧ��;��3vo�������ތH�G�VTP1[Ĵ���6��kƬ�/OV���fk9c��ٴT�L�����[q��]����>���H��E /���֑������0��#R�����Y6�L��F&Ug�L��q��t(AӉJ�v��Լϫy��u�gYX�/����Ĺ�kB�o��H�n��U�+��xҔC���Aa`t=������U/ʮ��!˵�ߟ���v+Ys���65�����q�-n��Hd�P�w[H�P����|��P����F���!�ۤ�f4�v��9� �`��8��]&�JzڭˬүW��ܧ]"��!$�1.'�K?�:�N�[3�&���ƿ�6.شd`��b1��DQ�4%$��{
��@�>�~W6:|�T��ӇҲ�%��?]S����f���`\0#�pWx��Ha*?2Ss��GFE�S�����r$��h��ܝBv��X;�yl>�T���"��O霵r�NR�4�QTcT�o�`#ew�#M�yiu�c!ĢMg��1�Z�)b���q@\[=)�t�K���J^g���k�8Q|K�XS��<'� L=4'}`�'��7R%>�����3r�&!]�3�c��s����u�����F=*����ʱ�@�$����2�k]�����J�@���]������S�K����u�q]-#Ut��_���k�RWp�km��vqT� u�!���{v��"_9:��o������D���J�0�{�X����T�'r�7�zb*�� "s�%��3����%�Gvx�]Ñ.1�F;.�_
r���'��w�~ �E;�iwLo��r�a ��V���]E����oD,-GTL�:'H��@�{��4��6��)�J�I�:^�]�<,���TP��~��k&��|��7��2�mP� ��R�ԬJil����u���q#m�J����}'1�7�wܭw��Sk`h�?�<�./�fJ�;Г/-f�Gt�UP��K��ӭH��a$�����f�o?�j�P���%(�Ϝ��R���3}N���NŷuG��l�X�)�+FwFD�]�iY�_;t��w~�y�S�$4�c:�]��9����eq|�A�V�����SKV����I�95���J��L�
of����eW���p��3�su2K�z��,�Y����uZ!�"���$�w_��[:����_��,�R�73>۱��(����ST�U��-�<N0�.�K~�:����*�:���&�!H���5�>��]���H�J�)e�i�|�_��}��[|��L|�.����M�����\��y;o����H��g�I�w��&	��v�CO��g���G���̮C����x8F�q~]��H/�m\�:�H��|`3��3�fB�xM�w7�C3}.jun=�I�q;>��5I�w��@����P��(-�J�2DZ�s�K�Q���9��ܩ�˿��zg�)&|Y��u�g���:�}&��B�&�T�'�K>Սϻ���\���a�2܉�2@�"o�
�6��cD������H��vE! ����#f��F���3MX o��5x2��|)���=v �F��Lm�?�;�LC)�p�0������4��)�����Z��%H��<�p��@��1~w��|�;���f��>90� ƣ%�� ^��cX����R�zw�y�l8B�h��+���k�9|o�wsl($J�պu��6H0j
��C�v�tP��c�B����+$$HE�-�ž����l�3D��x���RuM�x�.���P�&VR����6(�h��a��	f_�j�+��@�8��&(%b}�Ї�Q87�X�l��tsf�ˎ<���{��DeqTމa����y�����M2�tl�+A陁M��=g��[�G��G�e��7���O4g2�i9��{�6�С���iN_i�e�rv��#�����`*$sG�;��W���qb#\�Y��q*��9�mdr߉�o֮�0�� sɪyIX��-@y8�C��wi��wt`�h��-�u�w�z�Ӽ�&:�s��|�o��&�r99��#߁�K��(�Nֻc
;�@#b��?��U�Ƀ��$�-��961��"��C��Zb-p�!&�ew���+O�e��(�ȍ�xO��(��-���_\��[H/�~�O=���xc&:G� r0��!I�~�Oy���$v#q*;	d������#�����+��kc%�%$G2Lo���@m�Bh���� �Q�U>n�Y>#.�bR�qVW�:8v!��/)vTg�P��W�T��tB~������4���KZ�����j���s��*�����u�b�k�t37�����'�c돟������&d�Qc����o&�_Uh>�b���%W�|ג(��i[���#���	M.�p�[��r"+|��@�z'б���V�2Ŷ�R�oz�����U3`L#5K� J3��E��Hvze�G��0�A�ia�6�R�Q�������l9�"�� �\qD�c�����$�Y�~���*^~.�h
.C
� �F]FW;���L-�������A#�M�Nz1:�W���+~�E�l�hGJ�Р�Y����=��r��N����������*%ה蛢.�ݠu��ډ0��5E�����g�$	�[-�Z`sz�b�D�H\�������vȣ�I]'�6���gA�\�x����%Q�u~.�˟2�&i��Ef9�=��!�ѣW�0�o�6p��9�vR���O﯄`�4��E�5��㇇1�φ'*�� S�:����.��T[JA@p��<��g���'�W��8~�--Sc��?h���0��	���ꊥg�8᪅u�YX�����
i��oe���C7�A,��w�A;m���u�ϳ��zT��*�������a|�*��c�@��r��I͕aO=�D!v�y�!��P������T�Dϸ�����mf�NL�鷠�;C�{Ӣ�G5��U��x�d7�TD�#Q�6+�r^�˱\��꿓�E1�U9.��'c��$�j%�2�#ѥV��kz�KL��V��`��j�=��
d@��T�J6�&"�ƹCn�j�P�k� �;��1#u'�(�.���*�ˑ��3�ބ�G}a�{�^���wD@A�r�I�~,xY/
�����7�̅�?��ыv[mt����{���e1i�G'��w�n��V�B�J;Q/��r�YQ���u��V�
u�%Ŏ���F�Ol�= ��KB5iۛ8��ު�|�4~12����<j��t��8I���V7auU2̸��Ǒ�Y�mac�je� l�M��X��V&�ߕfl<Lj��j'q$27��ssx�/������;-Ar��:�)FEUt���J5�L����A��0��lf�o�׺?�VV��H�M�8>,��5V�K�������}���rH��鐅�o� \猽ɑ�*�"KӦ���X�����8�p�2�o�誫s�hj�ϟ�����1�����l��g�p�����k}�Ό^�Y�+�q�bky�̑�:鐲;b���<r2d�xo�I�og1�B!T��lg-%��8�?51�W�UM,�3�a������$����T�Le�^���IP�EQ�d7e��]�)���k�:X!����%���9��٠�ذ�g_G@�`L@�-\qR���_�c�U�.�l��IoU��X�D;se���䴰��ݺ�gSCfu<o�G��L�YL�@���z�$[��� YWx'Z�%��M�U�~�}�;��*	WV���τ0� fDRp�}l��%u��I���������a�{�#7����PH��Gz���5h#�@=縞Ŋ��_�����&����g�[
�O�A���0$��ߨñ��|�ǡY�
�Բ=�Nl����s��6�B�Gw��X�mn�M���O��7�
yՒ���_�zs�W�GX��g�9_ <�����3S����L���m�H�1.��DE�ǔ����W
�@�GΎ:>*#R� �� �_�I敘�dl���0��my��@����+q50�<
l�6@.�g�tis��7S���߽�XARl���5�4���٥�m*Lbh)��=]����������vs+�tX\d�Jv��K g������n����	��u�-��ҽ��x9>`�?�FDHS��P�>���2˴�
3a�R�O@T���/�s>`�ӪѬ�8I�V��(����q�)Y'!�?8��0�C���~�*w����u�sb�#��#����}-�a���Ûn�ͼ��n��F�������zE�/^؎�І~�1V=Ľ9T`�Vj{����m�%��ޜ��6���1R�l�7bu/�9���auBh�='1�0��AGg�b~�'^~[\���鐫��v��{�Ȉ�'�A�����v�-��f���(^8�э�͕�u;�2ˋX�K]^��[c��FS�M������� ��~�"Y`�N�C�<��-%F4C��g'c��� ��^�6���NN0Y�^kF������νlXq�����ID���a��MC��Ժ�� w���x� e��p8d,�/�`���]u!O�~=��\q9�!"�H�x����z�E<�"/)Q�D���O7,�>�ߊ����ә�2�'N�1���J��8κ	��{	��L��+�Ƽ�:�c�CK]�E��ό���H.���	H�H��8 ����#G]$���0|�zf� j���X�{�Z�I�-������]�Tnˇ�=%r�ōۥ����Ip�ё(eHj�T���}��x����N�f�Č<tp1x�b�ϭs���j+M�Ya�k��i��.�;�~ƪ3D^w��f��W(�ʑZ�
�g��' �ĖK'�K8I��	���E�.�kh�x
A9jr���L�c�ge�
ԅi��N�����ym��B���"�b��#n'� ʯ�#R��c�i53{	�
���̌���?i!kxa���H�8s����<K�d![Y�1~9e�4�ؑ�<��Q!�����\Ԥ@����u%����vO9S�Z��n)"�N�����U�	�(/�
��t���>ɇ���n9�w��`ChcZlXLY�Z%�6MП�[�����e`���nL�;#%�"l�O���飐�;���N&��QK`ԛ�;�����n�۴�TT�7T3�B���
0�C!�
����L�^�AQ]���
�UI[��F~΢��2/Q�g��#}���n�k���a��n���-P�O���j���8�B��\�l�!R��P����i>2z�����G%�co8�0�A��#�h�}C����+.E�9�;�o�5?xڿ���±e�#�9�e��Z��k7�0I)�k��D�,Z�q��عh����rƄ�#賟db;�k�n�)��������	r����fJ�&�&���*�vL�(gqOF�7��n����*����[γD��_+��Q��M��Ō�K^����ǣ4�!}�e�AT@��M�g!��g��CH��*���$� _���p�&�r�\�4Z
�!�p����azi��؆L��4����{*sf��+]Lş�X
P�#�H�ҩ��%�_fL�*���Ϯ@�1U���q�s�s�T]��-ru�-��K�j�xS+͠� 7�M�;dK�>N�ĬN��_~�lP�u�|<���jY�F��.�ͯ���xl�׃L_�z�T�a���ɇ�&��P.|�sfP�ݥnK41`}�V�֎Tf?�o@�� ߏ���Jv�01J�Ԃ�[C��[��wTY���<=:��������Krgh_���:�I�W���o���*'���rQ� #��Ԏs����cn]w���2{�dGTT3��y���b��YN�}�P|��88V��Zвڹ�0	�#����r�/C]l3�P�ɕ ob>�&���'��mW¡ǩ�W,��9}U�=�J��F]�!(��8����T���KX4]u��	s<̢8��U`)��"�)`U��Vf	�*�7z��
��=�Q%wGR���3�k�2XX��>��$�>dl�v��0z! ��o=k�\�b��|B�Z�#�Ⴂ�G��gE����/�����P- �H���೼�2p���3qLk%�ֽ���Rte��d5�p)e�V�T��H������m�o�0�����
�Ty���!�TO�rVX8��QpDR �ݨ�; ��D��tt���6~m�	�p��4P�-i�׀�ж�o%4���Y!���c��&���a����4E)Ϊo!&�K���e�E���fP�y����}��� ��G�D��������������_��o�M�5�=�1���f*��`��l���}�|,�Vvq
tQ�<ܐ�D���_F�w�!1iqz��28ps��F���@�y1��z	�����f���`G�t03�y�8�{b!#О�-��Ң`<铄�';�Ƨ�g�Ґ�1��	�"X�Ox���q����蚎.Ӳ�1�(�%ɠH�9��gz呤h%S!���u��0�k��0a"�~��N����^��'�cаE�I	d��7a7	���L�@�B}i� .<S,)�(\���i��5w�	R۔nM" >�#����Jkşaǃm?�G|(�l,���k�#�=sfeэݑ�#�R���傜�C�#*O�9BwA�܏����pAE���K�3�/���ǯ�o`����ܟ��"��u�����*�r#K���_�A'!���p�>\�"�#ˤ��w�GB��d��������GD���C�LQ7�Ll0v�q�D�n��&d[�ca+��I�VU��)����lo�6�����X�¿7�!,f���kC�yBy@�񓀢/�wgM������{<3jr��h�qg�0
��k���#Qt0u���9��Ř����Ż"��e\���V(�c�W�j5�L�����W��,�Sx�X_�M)�u��B<ug�p�y_��GW���)����2޳�F,� G��l�ƶ��<]�f�_�����ǣb�6h"L�@b�,百�#����8py���#�y��j�S=�Ї����kp@���Fs��@�T[S���aG��D�B�Bi�{��b��0�ݳK	�k���X�o:���u���/�S4����rS�fR�G�ɇI�v��6~r�峢e���a`0Q=��!��Oğ��4�ފ�USc^#�H-�pg�#���ʍ���k�$~��`uBQU�u��lJ7R�I��d�@�vV�����=�F�v/q��hqr��� bk�Ų���d���c����@���C��Ƨ�K�:M$3��f��n�G�e��QXa˃e֞���1/�A�29I*A�gi�o5���5_�W�l��65�C4A)�C�+"ĵ��8Y0sȔ���<��.j O��7o��bU�w%��J�Q�1��ϔ#�Ng�g�<���\\�R!�k�O&��,��GI�?��;��Ȝ Ōη��z+W���{X�O��U��>�o���#L�I�Q���p�ċ��~*����V΄mh�t߈����ձ���H+�[�P��շGN��1���Le��~�'��j��-�^B��a�f���P�����)���`9N�)f�6��k��z�f4t��1�;�^s�+�smj4����Z�8��Er�c]�����rt��l����uץ��[�nW����dFdld��G�C#6��q/~*�2U�����+
Ѥ�Z0#
���0���_�gM��cG���K�*�îm�����ml������"݌?�x�+GDͲ��aH���O��&,��VY�:&n���^4��d�����
����&�X�E҅��ˈ��;��ƻ�4�ӻ�@��m.��g��>:��6܉JkĶ_|�p9IC��ѡ�E�'
j���N~�a�
�o�QM��"Eڒ��b��lWp��P�G{*�:P��ؿL�9LթP���.a ����z��z �T`��A�i%ػ[�y762�(S�ԑm���0��h�3Βr���+�:��
�T|����U�*N�=^W ���[!6kU$m2\��G�|�D�#�
�ea���y M����P���1ux6_JS�:k�p�����ݸ�涚!Һe!Z��bd�0ܗ��]h�K0�:ڪ�-��+�l
�2&��e�o=�U�˟�ß%5=����Pt�4<��g�'�E���9{��=	L�R��ͯ�T�P�$:[ݫV�%�����Z����HJg�&���a�!�c�:�詪�n�|���o��L|��ɘ��/�_1+����w|�R_O�)��k^��	7�[L��$p$�,E
 �G#�J7I{��b+1Kݘ��$).}
���� �����6j��3muF�\󊨨#��]4[!g�D����x��<���%�Hզ�����KV���(��t��h.�������4p(M�`/��W����Yk�ew&��8�_�e3t%�B��F���������D�ָ��BQf�2åť3��ekR�roī�w���/"4Fwn~T����˜�z4�gZ.�
��D�_.��dZ�/C��V)����Y����:��C�æi�<\�0I�[���9�iz�.`�ve|�DH��!I��W`f�#�,�����dC�5A��+�����Y�-3L��Xʧ���jku�f�>�6A��d�4����e�j|�hCtSHHݓVU�O ��u17����7B��r[����৹���������%嶏_$[�$�Փ�L�ӡ!�R�(<QO���2F� `���0Ē��'|�Š�#��>����q�t^]��	�?��y�rkĨ�s&5�6�����/&�>�&˧��;B�B�:����g,a1���|v�~z^�l��'nY8���д�=	�f&���·�6�_�Wmܕ�8(t�;(�.�0/a��@�E�uG�V}�z@_< @
�_�9�D��_v�����j�S�.(Þ��2�Ʒm �64p�]��w����a���:0�6tJҪ�=�ڱp���U�����:��H���Ǔ�OUO�,k��F��D�8�|r�	f��5�c�3:��� l���8}{���w�|O �{7�g����U�W��8�UL��N��,���|�2��-��y�%M�6|:�W��Gh����T݈�[ ��,M����['!ɭ����@�����	����^ud�#fhWu�_���U�*����W��,6@��H0�:�]���)\����5�x�o4k��y�Z��=N�F�Zҫ���U�S�W����l�BԽy�E�}1u��qY{^j	R��5�Q��n�����������`o҉�ū�sj��pS�9e��%ȍ� N;_�9�U����^�F2�~��G�`g�9���:�/����S��$�=�l2y��I��&��v�B(U��dm1j����Q�c����C�qN?��]׭8�)%Xj�u~���&�S�������q�ό�w�����.cR�y܄���� �#o\����D�/�X��'���*%�UZ�-�+�[��څp�M�⿖.��6T�)��<�\qZ��|���
4��s+����)P8D��<��³Zg����0��x.t�'CrꚊ�-��Q+b�Es���=h������1YI�~��n�3n����°$u�.�5�h��1��f�r�����/F;p�L�$'a?��t��E�F���~'�=�(.�����\�,�����E�S��;΄����F��>f=�(��,��b���C�ڄfҍˉ}),�n���qqqv,�7��շz�i������#9��k��RC�!�G%P�]	�ę;Q*���c�HB�)?e�՟l����c��Y��>���q�6���w��v U�USlS1��	��`~��PJ��0���_����m D��iQ$��ث��ۉa��Y���(R��ag�{^�g�vM�Z�by\@�CEہ�(�<�����:[��Yct��̀,���[���d��1�P�Q|L���-�~���0J���+����֨ܧu'��F)��@�����{EBn�Ķ� AUE�xM�\���F\�!�I�*�U�^�������ۙ�����������JOL�|���L�(�u�nm��Tܣ��[Q���$-�&(�|���{/VY�z�|w�g�*Q��V�t��wU���Ԝ�xw�������� ow�hG��y��gZz�H��ry�;�_�n�f�Y^��Ey�Ҁ]'e�I��*˜���ml�0��VOm��_ �_��w�hf;�\c a�C~��b��R�_�j�Za��Zb��i�� �td��3xZL�L؏��@��F�4TQ��i7��dh�jfh��Ԟ0���e<m��|�]���ʴ� p�W���(!�D�_J�&Ǥ�rI{n_��>3 o����~�\���W�M�O<��Pl���[\b� �~����mق{T�pUp�;#a[�(3B�wx���gV���qʖPH�R{*�
J�Y#b����H�P3����I�ZW>^MVf����$%��!����^Z��@5?G�/�	�۞}V�=��0�0��R�"*�.��Kb�ְV� �}�8h&�z�aUKyc��`�!�ށ`�;\>A�>UC~x]M�2�����5_:��o'~}�ِג�E#V�@Ԋ/�T`5�B�^2�����fs�<pEj�?� ]���͎:��rʟw�'(`���$�5=��/�<x���UJSƋ*��SI�L�T|}�}��r�ilѺ��K�\�,9 �~��GR ��Ʋn��},�~FP����ȭ~p��Wk�����1n�"��A	���c�'b�{.�'�x���n��gK�A��.�����D}�!H����nE�ɐ��B�� �]_!o�P��2c] )6Y���*���F�� �j%����}s+SbA��,`��(�|
���|���LΚ$Fej>Z=��N���פ�
7on̒e�I�i�F�׵賂H:�ƕ�a1�oY���)�-�a�5���d�J9�2El�fuj����|9y�^5R�":�z�X��<\�~~��'WʡS�EW�r��1�0R8=�9C�/�$ϫ3�{�*�`͞vՅ+�Z��N�W68�F��i-�?��b�L~�~�^+��>rGߨ�Z���brp��@�&b��NN�_��m�_��s&���X]�;�;p��|�B�6]�0�3S�@.��3I���9��" ��P"�]��K��m)5�y���X��X;6gT��0������k�\Sע�/Q��I ^Թ,��ӥ��jrOl����� j!���D�-�qM�^��֡pAp����"�b̽F�X�p�����doP6_�M����4/��c	���;��*
 �fh0J >����W�y��+�E��������Q��"��4%?	C����{�L7���U'���܊Qn��v�G�$f��ׂ^����l�C�x�^�S&����֖�Wß#��V!&O�	ʤn�y�ZN��'Bm\;q�0Q5������E�g<j*�~��䁱��r䐅��צ��Q��nbj�q��FLw�r�2ګd,4Kn
��Q���U@�>FZ�N�B�?M�$D~=0􊜦�.F��+J}���wEq�^�-l}�[�ۛ_��ǔ�9�f]�1O>.�hd�-��L�W���7N��T<Y���ٖm��G�I1����	{�Y��x�A��?9��SZ>�@]����BT���^w2���E��܇B�K�x8K�9͐��2b��h%lR����<���e���c�QES�#系�C(]M~4o~�ʿAQ���N�U����� w�����>z�T�����wi���ב���r{�VK�n��c���:��]�.��[�}栄�����m������t�
t���^�\���z'�Z� ���ZP�D���M�T���2|~�2������ف��=T��N�6� ��J2�n���!�E�X�4�ĵ���3!C��ZJV;�z̺�t�y�is�%U�_ڑ��p�PRR�L���|��b,y�_�ܪ��u=�+�RQ��vl[�O�U�#��5���!jǅ�s�T��or'>ݱ{���#�U����v����7��q���4��X.,�,G�$�-3�wG��N	��9��\��E��.˵1*�<h5P�C+��HB�>�^�k�r�Ri���I�pqy��]�Yyk�j�p��a��3_uI��p��<��/NXEY�,�m�z5L����I�������)hq(\�L�L����~x����%�xwzD	�0.��0q�[c�DKRn4y�Y���E_��S���n�V�Z˺���Ι�L�Yz���?/�4�y��UwϦ�ԟ���X�|Su[\�w��yЋ��p	�q�^���e��k%ǣԁ#Er�(�bO�F�RR�]2}6[���`�WnY�����p�X�S(��51;����;:��|�.�Gh��&Q*z#p�U�3R횁N4��}�l�B^��F� Y �If��q���l�:Y܀���F����&Y#̔z~9��K��0W�ވ��ᦨ��B�+p?�����×�$����8{�W������/�}��s-��\���aA�w�*�t=CLY�+�x�)얼j�
�$j\�D��9����S�����1,�\��{�%f�����<:�%�325�=w��s`��^�����nr�JQr\g�5��=��>�Y;�il�����8�i�ύ]�Ƹi��K(�$��tX�|�b�wF���E�'��g�U�%�� 2Sp����}HDk&"}�#"Ņ�y�R{	@u�Cܦ3��v@ߌὼ6nt�iڐ��h��5�)�FwsY2G���B�h\Պ��6�[�|��G�:��kP1r��%������{p�����n�_6���h[Ջ-������z�6����L��T[��c@�:KU
3��bh�J}t�W>m]�y�-z�l`~��۪�$��fl��?�w����bL�Т.rL^�j�"�vzC�a��n�N��=�m$��Y�l�Fu]VFt�oϺjLl��v�%<�/u{ɣ�����iRT�=�	���V��!#ģ�E;z�o�.mΩ�q�M���礲,��e� ��G������OG��M�08#�Ws^����5v	ab�׃N�\;�Pqr�1�z@��1��ŴԚ�>0�~>����߶�j�cMd�����q��Pp�}'�h7由K�W� 8��F����ʾ����M1�ye�̚�Ϣ�SQ�q�n˙�V��B2t��"h�\�>j�6�O����c\QA��M>3��u�n�<Q���Uʉ�?g�F� �e�M����󅾊̕7H�ϩKX�µ�R�p��u"pB�=��f~P0x뜠j6��~)�,������p�����.�G3�����u�[9��o�[������Ζ�=���c{2J����>�Z����u���H��b3��F�g(뗊�����L8J���r�n�v���\�'6z3
��'
�� �E�t爘�yrD�N�z����P�I��@�	Bt`�.ݓK�镹�[��-�(o����N��z�rȇ���22��4vA�)���Zd�@+�-�����E�I��5`�}7N	��	��U!d���J���n&�����{��s�+ՁY�bB���/��h�z�s1�拪��kUܨ�B{k@*dZ�*��f�-�!�U�=�i��ɚ��L����u1�W&�:}�:
���Z3ܡQ�N~�	��sr����Xmu`�Jב�!S���N��^;ƺa�s�#_����O�{�4n���vW��)����x�8 �t  >�����wo1��N��zH�]�Jc�d:쵺����H����r�x����|4�I�\l�0¿ �Y���
e������b8;�[�D�
C�;SqN�-?�W5�r&�X��i1�[r3x����m�ē�aTG�7�B���3w�)�=b�qҿ�,��c�����4P�@�{[9F��M�{��^,���\�q_���Z>͎����`F��h�vҒ'a1qZ�\�p�RE9�����S�W.��e%2�yS�9ON��//�Nٓ�5�����ȥ�&jb��(����CO)�hc8�2��;Q]�^�59?u�	 �v�4r���~ڝ�����A'*�����IQ�K��\��iw
��&JW��z�γQ�X©.����O棸4�H��4��=�UH߮v:$���^=���-���jv�E���w��N�kj�
����=ѫ�.B�C�	/*��=���U6Qlzz��j���Ԝ���F�J`"�H�<������!��`����؈S�"N1��U�{m�����l��߆=���P[׍�_j��R�g�^~����#�,*M��1�߫�&{b�RץZᣯo��ă���H �����$	��J��t%j�Fm��ŋ�'�8��Uc&7�o����nmx��^��S������5y�,a.����W��x����yE����Y�Y�.�E��^��C��%2�rn�Cɇ��aC�@�V=_�?U9<~�h�t�����@����u�ak{�������i��˛w�j��
�07���:���Gm\�:��?Y���a1�`��[����Vuu���c�i��Z�f�'�d^&h&�,��Iڔ\�|���ʔ���T�W��0=)dut�g������4���?=`^���7- �>G}���^�	B�<��c��-$Y��f�f�t@�\���m2s;'�N+����]	�X��z7
/��!\Y՚���ܢ���Q�ʖax��{Jw�h��`At�� ma�\ �47�\ͫ��hg������
�)��+y���u;�+'�xE�GΊ�A�,��x�WL��8��W�d���TE�3�ݿf��f�c����
Y�T��C��w�7��_A��O�\e/��GF&�T9��)�Tꍃ��B7��s�J�EZ]瀖�y���9�%:ѹ��O�Ɉ=�[��`�щ�.Q�a�AI�G�G�x���ѓ-M䰺��a��K(q"��x�_�,�뢟��E'���i��N��R�oL�71�6jF��d���\QP�J�z� �,q��јt�8!
����Ѣ&�[a�w�M�r��ú.�I��v��jc2�\>�$���@���h��4��J�.�Nn��T���(�+�O�����|�L
ly5���j"R���K��ۚH�"�j�<l���&���Sd����������x3�����%*����B��)�xs���C��Rz�1]:�O�ft�z4���Jˠr����kNvP��E�6A�Kk*D�l����͌�˷H(�WK��j6�����Xڨ~�=�����ĥ�/ o����s����Wa��Bt#u<Z���O���-�rŊ1U�N ԉz]9Xg_b��NĵhA�B�4ɨ�	��C,�7����ꎤ�5Y�<���<�c}��/���Ɯ}ae�m��Qm��3����[��?��_�$Q5E��Z��)�-nG�AR`ҽE'r�D1�z� ��Y�Y���w����p �0��V�VKI����u8�K����Is���hn���o9^��z��֠[� L�`��|�
3�B���Lx�'�<�#S{�&�4��NʵR�'ʹ%���W��#���.�eܶ��L|�p�tY|����`�0GƱ�p%�k�.�ŊV�rq ��|a�zBl9�NH�}0TtK��fט>�&��U9�j�ٚ�5�U����2�.���L=�7N^�ּN�Xc_-�s�gz�X�Ybu�/��:P�a��	�S��\im1gW���^X%s��O�P��E��a6���BvL!�6B%�r��Z�`��T� �~�a+c��j��[d�m����UIb��z]�=ͣ�����|
9O�{��\3�Z6�j.G W�����-��ÝX�L2����GV��:1�\;��Ƶ�QZ_8[M�,&Z��j��SO�\;5��n��a�u�e�����Ք���c8�|��G���i�8s��Z �bL����q:�Ȏ��y��L��g{�riځ�Q��$���n>��Xk�y�"��/|3�y_yо�P���S���Βd�ýp�D�Sp|	z�f0Pv��>��:�߂��<^$�*��o`휏�z�yx3�f�ֳ~ bO�2��.JM}���b�ì6$̃^.���zң��i7��.���S՜���OO6M����|`��u��MV[�僆=|���|2<|^#Q'场[[tH�R���:��5��	��9�i}n����B��E�J,3� �|^��2#N�a��'?�5�j@�M�9u����Pu�������^��h�����2 �0 Sk�+$���_"� 8���%�����͹�g�c�k�b�WzZ�*��j5���6���N�1~G~U�ߕ'��JJv�aCc
�P��v�>�K��鐚5�
��#�Cq�/�<������-6�Z�*"r0i���a*���4�oW�P���z��=�{N�:ߝ��������Y��bo�^?�c�PxR�Rҝ?]��<S���s�/VJ�	�~Ș0'�s��wU?@������p��'��Tj�^��~���2��/h��p���_	�&k@a��U�H�d�ə�|J��R�vU����D��$R�׿���sX[->��Z}�B�\��bXca0 Y8�Q�>�$�zX;>��5��׆��2�%!�m�%�;��W�}:���/l[5���<v��K��s�kQ
=Oc�}�O����켤��#�����6%��V|yY�)U��L���Z{�Pi�1Q�1�w�S�k��&r�U4Bd���i?o��ʤ��������s&%�;�l?;�S7 �W�9\����F�6Yw5ݲ^s%�_�s�L�ow�v��BU����v�ʎ��Gk���%�T|�z���
���� �s��=�`u;�@��B���C�xR)y��g��#�,� Ģ7�.�ˉ��{ -�Yل��T7����}�!�YB�o�̂�bMi�d�t ��  �9U{�E|�Z�>,L��D��� �ݛ�@�����F� ������^�LR}hKO�8�F�d� �
��%�h���'�
,��{�S٢�x��#���BO�\6K��^k��i6�t�ja�P^，��v %l�i�dv/ʋɱ�����������EM�J����Y�p/O~nŬ-�դ���iNa�#��:�j	wyX8cq��M5���l�25?˷�p��nY5p�����T���H�՗�!�1�9$9=6>�co�kg�0�����=t���I����m�MU�]������b��l��s��٩����s�׉E�Q��F�h�|�T>��a.����}�����A�����p}}E�Ω�{_�	+��spi	�I���}o.  ��	AK��>F�@�J`\"=d�y����+g��;1�Is��Ű���@��:BMgK���-�G���
�6�&����)����B�*	��ŭN0���lw��I/�G�ЪM���H���~���?��B0�����o .@�6�U�B�{�X2�8p��1-5�7T@���
,�����c(��H�艎i)g��%DddI׹>���|t�b�ý�#N�D��̠�������x'�B�TF'k�byտ"�^�J�ĭ3]^a�&,C�+M]���S��!wRVHQ�>����olj��w��F*������_��3n��'�<��a{��D��{�L-�W^�H�O_�#���ۜ($ +�F��}b���p��NM���j%��P�@�Zw�łw�wSG�*�#0*���'n/�>��=��|'D.�e{奠?/v��2b�q���M�7�ט@���HH^g�i]q��*�Ù��k�A�2f�@�0Jm� Tрۣ@@����)4���r�' ֈ��e��LZ�G��u�1�Ɍi�!?Ӕ ��mI�*�j�����#^�oC�K�J�������`szy�,Џ�d�N�"���㯝��"��^��m�u�5�-� �Tx�b�ߴ�u��۝�/���2O����+�J;����6�c�&�`nϾ�%����C�晴�����߹����̢�k��h*~�xQ4��l|,I�c����R��*�f[�sޘ�����E�afG��J%DM��d~0�ߢy<�*��$*��cH~]<��rls��9k{�u�d�6��MY�C`F/+���y�k2�vW6񛓚�g�Mn8��� ����䤹��x֩�Rѕ�����=O�q8<���J}�pJ���W�X��r.�za�ҿ�8�������#��s������@�gm���`M`�h�����V;�8��ӷ�o��E�^	8���I!�~��ks`[���u�)�m��ሜ����,A_�U�{4i�z�����AkA�"l��tf#�VΙh��Z.s��@E�zS���OҮ��C��I��\3r4��'5Q}��&�=f��k��1ȼCn0̘�<%�t�]Bo@A>�u4�/xa��ҍ���2�V���]��d��[>���0���,Q��Z|9��~E��܋�B���MxSSL_��j �|[�����"Mt��F2��_�ƥ9�є8W���A�����@�ۅ{��&��$E��f��jRP�K ���݂�3Һ��t#N���֍z��h�sO��t�a�K-���o�����@T!�q�q���jx��k�~Z�'j#N@<�{ߜ��`��v	4�	���O��i5����R��\w�5:��5��ϳC���g�YE+�������@*����c��m�8[-;�0"9�c�n��/�ܱ�0
{�8�	���g�B��!�x�]����	rG���
�c���g��Sk���
3�ZZ'P$�эZ>���&�L�����ʝ�t�J�Qs_�~-�2E���3����S��_��a@�<>����s^G��H k������7��s�df��hT�l�H
a��|l��y�@�Z[*�e*�T7\WX�ц��+Thy)�*bb�ȟl}� �Wr�+f�mRn�hr��I2| iO|�����y��{V��7P��3��������0�#N�|���c��!n�5����;��ѳ�uF���Ƶ�f��:�K�"�lp���dQߤ� 2!�ij�sL�!��f����2��H0,�!��?QFw�.M)�ေ�d��@�VH��h��]3(�{�ͥ�?�A�`x$�qo�V�ZE��+0�'� <�j�
h�'�dN\!1gs`���o��Z��k� �>Q�_��T��'�G���>�e�k>R!*o�Zu�P��nfq����	��Xî��G	�;QY��)Vr�6�RdN�Ov���4ւH�rq�,���e��j��X6L!�>���*Q�����2!�k�����6V9�|V�c(���?�L�,��9�
klG��"�yJ���+x��y��(�V��aȮ��-�����)lE��u6�^��\{G�8mNTB��U�[�.m(SU۾1Vk1�j��̑��<,ۂ���pDd�]B�E1�ci�E�@,��kJ��\�hI�b���$+>3I]R�o�m�Ō4���$�|6�nv	��F�>�+A~ƚ@QQ5DOl�&#7 ��/��Lkȩܢ���Ko�]�*Q���K�Ϫ�
���P��i*%7��F��A��0~"��w�w��b>�\�bD���:ȯ�&t�7�g���idO���]kM��G������5 ߴ�:D�K:y��z>H)mm<}+AA��6K�������1�VD��-�A�.�%%�s�cz��!�d���5#��j������L�q?F�������t
op�R�J����c���G��ύ��?��/7�=L�h�E�)�~��U�,�n�|�S��[T������J/�QR�Q',FztI(s�����,����I57
9z��2$	��W��$~J/Zl�_T�dd�Hñ{�xa�!��w�W�?;�!<QxD�iv��ڃ~]&KU�y=r���O����v�㙜������c�Y���*�-{H���� ��Qz�r�p��f���$˳bQ��&��`y߂�R��u����6a9q�W/O�����qqd[�I��s�#��a��i��RC,����%�[���آ���3f���#���tE��:?.1H��a��`pjOjګ}�p��^*ؽ � c������܄P����d�jF�v�C����Ok������6��:�9,ٙ��_氠��x(1�����-Cg/�}����rj��Ӓ� �_U�� ��-V��ʓg#��[����Fj}b�����s<��J��_ٔ�D$D����nv��S�v��i�f�.~n۹{���3��$�PE�/�2���%>��뮚d��Ǫ^��(����,NPT�'�c�q�A��y�c��B��uw>#|�-�A�H1��e���aq�!����n�i[��T�M�5���=%GN�abo�(-��x��^v����X)�`�~�\K�AG
��khif��X����{��p��lh�Dʑ�22������)�%��9�������i�.���y/�Z�5�xu�.Q�_�'��
6�I�pk;	���Fs�S�[�Ҹb#��z�g�ygB���l�����/�d��\p�P�j�{Y�GN+c�J�� ����+�����ĠQ(��zb�<kB'o���cZ*R�r���8x���ds�	盆�P��yo��Rq��O8�ֆ2_ò�s�C@HY��E��e�L�7x�ԗ��u�C"����G1U�#������ҡ�m�0�iBa���o[c���jL�]��k��g:=�N��r,��Z�1���[�ݷ;�)�l�Ad/��|�L�&��8R�B��8�_g�"�w�#S�Ќ��dد�v�kl�K�z]2�X1�4���}q�XA7��]\O��`��X��zv�&�^��6Ղ>��
T��]10W���>ڣ�'@�#��0��~=l���g�m���gFmV�{��9�sKtU��?��8�b!e4�X�������S�pk����,WI��~�Z2<,z\Be!S40��(y �X�@A%�˺ڰ��+I>�4����C�秝P�G�A*Q�L>ȉ�����dhF�|��E<
Λ}��_-�ku;%�5xi�!�gl�zL2�Y�5�$�>Y�o���\�/�M����8q���ھ).Q��nQp�z3����thޏ�͹�`��	�Up��'g	���R`1 �� o�H7�1��s@��ƳE-��dw�ACJ�Y�
/w2���_�8e0���8�ē��O m�o*H3��L���zw�dQL����Դ3nh�歍?Z��_�� poH��˗B��<Dnq���L2��9�ʬ^)q6����GCL����5�;���Y��V��ְih���˸�b�v�0]���_`ԍQ�S��L�fM	��>4.�r��?0��~����)���V4	uʉ�"���-������fi6,
A���z�&b�o�^.��T�1�駐�`��߈��O�@�����Ly���b�qZL��}���˧��ۑ���v#�¨b�:/�L��=����u{x,¹��kL�����(����}�
�ɘ!�V�@u�5�Ij�_K;���=�i�	E�-�v�>sᴉx�����N�{�#�M��F�~���a1n�*��ܲ ��[p>�>��ӧ�#:CDA�9 ��_K*�I�Kw��Z�>��/�рC��VY�mC DQ�f�T(�*&f��~��ڗ�ڜ�C�6���e����(�xT"O�����M� �TG���JԵ|mt{�ϊ�=�Ã��EXBw�pZ�ؾ�� g������&ħ���RY	�$F)��F":w�Ho�m�U�*����(�.�P�Hja�!!�" w��%@���	PT|rMG���z�+��ldbo�����.*~O</r��� �q^t*���g_�v�'��]�+����6�$=�;$ǻ^B����C����� ���GN��O�cD�V�j��ϗ��X'�7~?�\�oY��)x�	�e��"��u+ؒ��g�,&��N�7�J}���e��K�j:S�J���cE��o���]��<���8�Ou���	a�����v������蚥�{wQ�qo_�X �{vdW�﷾���~U�;��@!k�헌"�mC0���B	������ν�o���:!�/	Z�h�/x�?-�e�s�U�x��c�C�5��c���!�z�L5�s&I�#���Ai��Lw8~�X�!����_x�����~2�`@9���� F-��k$��ھ��P	(5raH���P���\�b9���J�m�5��H]�pbr͠�Q����ο��B�g�����rkM���e���SjT�:���� ��AȳC�@�U7���� O7�Qk|�2�U�򄁰��,�LM�F��M��*4+�%\�y/�v����=�Hcn>�R�)���8}\���#��)��F�`j�n�
3��������%E� �z4E��S����a�{�����:o�I�Ѥ�K���Y�^7�`��y���=��=�h��\�[l��%i;��.L��x�Zmwx�sx��)���[|K���E�K�.�����c���v�\�ӻ�@���}�Ud�7.��4CᤨM�.4�l֤0t�K�$����y�f]��}"萒��y���W� T�a�"=���a�e�x���ls�Ŝ��U��j�	i�3�Y�}��A����I@:�=��ש�v*�gPI�����pIZ<ݭ�"��%��S)}�tBe#����w��@�1�41��|>�ߜU��ް�w=P5�#'N���ϙ,6AI�B�A��-�����,Rb-aWl\y<��N/�/�<���ߏ�^`�� I����
���yڐ��""�tW�K)5h�+))���@Nj�x:���Ml%,K$X�$,τ(�s�U����g8�'{Q�یc'��¸կ8���N^��!�y����z�_��$\hi��(��<a��.�[%P�
�̴��vm���x@����L��D��a {��W]�j��� ���_��~Y�r�W_�r���*�^~�'Pɗq��X����V�v.L�_����ϐ��%��)�a�~����+�p��F����d�p���f��@7�R�AIO�������}��F^t���P�M+4fm�����x�䥊��p��Q!-ON$���~��������G�cV���.Ӽ�sQz%qV��ʫgv���ѥ��}��u��z�m����� 췬B0jPy���S�U�c"�	�9�ׁ�.y�ǎ���2�G�'��e�܀3S6p,6k��S"CsX���Z�٦Joͻи�'q89A����x�<|8e�)�k�	$U-aO�������jO�h#�K^������f�
���qF���-I$ҩ� ��~6��CݚV�ݳn�2�����-��^.*����'p�}���%膂sV#h5g\ȕ�)�N�����챇O�D
����5�l���}8+O+P��7��:�]E,���Zm�`�,�.TGX�q�FC�I��̾i$�Hj���|�����
���8Oj !�s��dՃ�f��"�|OƑk��U'ߥ���y!5��%x�d*��B~\���¡E�ԣ��/Lw,3d�;Hс��i�̓2���;z���Վ���}����(�w7E|���t����w���~}G-�l���X���l4������z���-w��L�B�Z��{Cy�����߈���~�9�{@FMs���h�*�z�%�J��KHIn}��eh0�;pv�a0}4C����q	ұ��Y�y?N ��N!�d{6{,��q,�6��X�]��Bf�9��d�����h�Dx�2�������䭴���dL
��a�!ɯn�����ٌ��ݩ O|���u��o�v����<�2�>/�<����V�c��&�`̀C���[�������ԛ��#�Z�O}g� M�����]H�u�x�o���+E���uO�)^�Ĝ$�� dh�DE�讚�|����n�g�U�ho�+#�>�ė'j�|�cdj�q�ĭ��U�(˒~v=AK5d�z�~>�z	7�V�kQ�(N.��Ic"���7��
�v�Y�Ȃ����@���`�z6�',C���u�HܸRv�l�s�h�Hp��rE[�ekdN���f���"bB'R:��1��ZF��^,�%��P2���m�FQ%R��t� �I����A���u�瀎,��'��Q�1���<������`9Nz�8��%h�}!llH�1κ%
O5q�z�c}e�}�T�M��j�^F`r�{����9�����õ�m >$��'�V� ���O�U�s�(��R�)�I_V���&U�@�M�j6�a¯a����;7Ǯ�^EƉ�+��cTI�4"���꘩��]LZV5{U���
z�]q�	���i�݄(�OJE��&<�^ �#?{W�'�F�T�vmgf5�����ƒ���M�6pI�eN��š�X[-����~������XjwKkعt(sub�~������&<&��Ka���s�P��b-9*c6����wP7�;y�i�	��S�6e�#H��b��?/�)P� }8�(����jz����m5�	\g]t��4-p2޽N���-'g�<eU�j��?�H��,]��#�u�5�#Z�Q��+��kJ�qN�}����R|-��I2�ʦ�Hڒ��&j�y12��I�q@��	����5����5l��4����)�P]�e���t�%�iK��2Kox6��OЕ,�-S����t��7�����?"��qVL�l/�S�%��������#�-FH�Q"��)ȝ��:��p��.�#��,���x���;Z��3�YOI��� �v�uR���Q�_}�������.���[�AZ[K,6J�5 G$�v��?[ȁ�+��h���$h����a�`Y"����Cz��u:��]~����K��Y����!_�ੂ�����=/u{�	5>PTI:��bN�\�b����㏍����I����F�>�ŝ�EPa�aܿ�U$��bp@�*Q�e�N�+���Z4Dߺ�Hj�>]�"��g�'��  s��Ɖ�9�A�W{b�յ�@���a|�
p:<�k����P�=[���{�|���,hƀ��Ǖg^�l&�u��JJ�ہ���A���O�x�8���F�`�5z�>�7�_{���ӝF��F���b�s�)'�}��JoQS^{ڲ���Q1������EY$�K~o�M��KR�9�B��	ް�6Z
^_^mCE�
)��(�c<��!Z��j^i����c胏�!�#a ��Yo@�S$X^����#�e���Iׇԧ�ELxTE��3���h��1?2�>� t�CV`�X1c��+�����X��߰�P}�Xm'{;�!Y�>�jH�˟oTm���f�xӷ���*�:���ǳ�"�@4M�،J�_:�x���Q �\`a}������
9_nV��!>�EjW�mD��O�v�%�ǂ�О�:���L/�}rDW���#D����n�5����lZ��+�ɪR�S59Q_\��	��/Y|&^�,�z5��6�B�QG-�z�=$�s_��6?6n���O�*�v��Yi���\�Q� o}�i��x#(�W���t�	��ã�*9^`*%����H�q	Ȱc��z帬.H�9��Xz��W�v<��"o ����*k�ڛA�EF�|�2�߶o<tS-�yN#���Q9��9���zȦH���=ͺ�m�Ȣɵ���g.I�bK���ņ�ԃ�)�[B�,3�J�
�%,\2YD*�M�gb��Na3������0��&�Ŏ�G�*}U��8�&�=��#>;t<���q��3�R��c� p-O�	;o�'�z����jx���,�� �q�y��uE����3�K(�$����<�~��%nX?�t���DQN'���K�.��Ɠ�]!�} ���no(�X�2}��zP��p��=o�;��,e�;���Dt�q,qDs@Ü�}b���[��Ű���,0��~ �	���z��~K�v�<J�	3ܻ�X�{����*:�{���PNU�0|k@��܊���h1���IIukV�vdS(�l�c�����Z˰��G~�]~ئ��ah-}�'���U����Kf�I�]�
��'n�\f�٭��|�9�փZz&��g�&Y�N�k��K���TM��},��Q �!pC�V�L��� ��/Yfk��O$��<0
%w5Si���C��|��K�)�ru3eRF����ߗ�@��ho ;~v2�I	,?��3�4��_tse=��l�{\�Y��g����Q�v�Z��� q�/2�Wr��.�Бg5M�pͯ�����++7ܨ0�lP�t�[�z�~�ȅ�0��CZ�	�F������0���S�"��A�u�d���?B�86U���g����$,4I �W���{Il��|n�XM�w�6�������	�k��	uJkq\�A�FЌ�b/J�Ｏvv/�%�>��5/	ɻ���3ļ���QfX����u�� s�%9D��}׵�3|ʝ����Ĕ�H��E��W;�ϕɶo�Uc���1�t��@����/�\2����L�����60-RU0,�����ϖ��|?��n`Z򺅩N��u*Tۻ.	�ќ-oCI���d�UȰ+Y*���ݹ�&y!�|ט�	j��i�z$�{۠yK�~��ڂ��;u?�taޛa�6;�S�荛Q�I0p�?H��dQ�{޽u����-�{v�L��9��W`B]��ynԽQ��l8E��0���F��wW:^3����H���.'4\\.��^FX�=95�0��c-3�(�x���mO���p�����o �^�20O���,��}�R,�G���c�O(� �>�!F�g��9Ie�1��+^U�k�m;F�6���{���T��@���iNFr2a��s��R��qf�+u&UZ0����sG������]th�o��i�m�~�,��&�m����	�e����ҁ�&z3���>3t���h���t�^�k���bH{j+���FGBG-�@nnr�����u�?�7cz�/_��hO k��������{�Q���R�6���$Z�����F�UFcw�����N��ҟ8�3���7��c;>Oa7��5�'6�����s��iL��[_K��1?�n��SKґ'��?oXU�lR
�Y󴸏VD-�"����S��?�/�e��4T@D�A�՛��|fh�"GR�`m��L\�~豐�����+�T&H0�֊X�������F����^��63�nKYD�h�t┉�R=ap'Uo�(2S}���G�-�O��V�x�����>����Y��h�H+Pc���V�u5U[� x,PH�9|�`~���[/����u��?��+|X��1r��c"f%Z�H�K�c���[<������IM�~E1�0&�)Ce�C�3%2\�.�~.6�11�]��.3�"a��*H�W� .����|��8�W�ʜ:�ku)� ��$�bo��:"�G��P���I��\�'>�ѓ�H݄�_���L�w�C�xp��1�4+�̘�t���0��@X�����N��Sz���#T�'	�x/�10�Qcb��)�8-�i�^<XR2wP��.���߆�L!��ī��MT�$�����Zݛ��ɓ�ŉ�>�M1`(([�w�G� 7�Khh��_!O}��$�0k�afī�ȗaq�=��D,��AR6� ��{H��2�h]�&	�C����E���3��u���"�D�M��2�%p���z�r>��`��R��@�c��a�JZ��欚�(KV"L�isC����b��A9c��Ej<2�6�N�vn���r)U���B_�����[���Q�w��,�l���U/��2�b�W<�7$;����B�a :I6sv}$'��� ��`V;C��W�C �O��_��ť3��wQ�g�`q3�_x�':�qw�/:yr���o�^����e��ywMI�����U�{���XsR��<޷�3���T@��� �~��#L�����}f������"�?��1)���{6��u��!3=�w&[ؔ�>?»*��7n�Lv6�]��Glc^���y���U<u�����9)��6%�e)�$��]I��*�Yfj �A���c둛9�Ҥo�ET7���,�	����� ����� �_:� �����3-���g�������9����Sz\���ha/�X�!�w�l'���� Qk�m���#%3j�j�5�";��L��Q�����v�s�d��[��ݺ�+̯��PV6�6���[M� \i�,���KEU��u)а�{1[��1yY;aD~�����S���
��jj0�}�C�������=������������L1���u~�9vgU'�'���"T�컯Z�M��9'� (N&xK� &�� c��L�a�z�lj7f4d�l�O&/D�(����כK�)#�h7�Z��e��nYǞ����-���r�J�B���F���~�Q�v̈́\��M�gP����m$���@�ӛ���O�P�� �ci!NB�����T���Z3���П�(e����4���2�p��T|ZI���49�z�6.|%�	������2���\8�ɢ�h=P��;��Q��@����B��!���Dpn5�u���yM�G�bc�_���H�3�1X����,#�~F Ė|N���� �`X��f���J�f�?��D�ƈ�",�w�8�G �f��Zn8>�W�b�8΋�}� v��������e�:n�P�����Zʠ2�P:��)�b�L/�&��^������Vi�<ɝ7�_��Gp4�4�M��kDEk�Ɇd��j�J^�����A����^[�~��n��$����� �r��G�
�$6��$����E��������h�m"��<�8��P��%��LW�7y�a����ҝ�|+��s�!�������b%�EX��T�����	+�J�$��r0A%>�쎑�n���9T\����w��Slhk��@q,q0�C�煑C3U�0`R=�2?��]H_:O�Q�YX�C�w� /]f�X���G@��ݹ�����i8:Xb�A@uD#�E���L[��I�E$��UE���h���B�%ᔪ®��~��c�=S.��/���"��7	+����5�s����w��f���T+��Z�^z7+Q����F�2d2ɲh�K<7�e�?8X��ɟ�	X�Z�a���V�t�������Z�|�G�/z�A+�4=���*�m���eYx�$�&ݻ�*����GV�1�������)����qS=�����5"CcpI.���B�4�Θ��ĉ� _��A��c�Q:C�z�M7{���{��t4W0Y��2hu%Gif�L0羗�{��x��p#�}����t-�
��o�&�ff*N֚���[���b�2����.t����V�r���S�����_��Aa�l5�s��l�@���8�n.�GQ��rB�v�q=#؂4���s
�J��	��o�K塩 *����Gl�6��*�e�7[��:����N���|�P~�	sP�t@��<���H�y{XҲ�怹��DS|�_�#idv���Ë&X(����y��R��֌��/ݸӤfwb�
G����2�r���PW2�������3�l�L4w,��,	}'et�z�ߪ��c�*N�������(���D ��*��U�����(�$Fi;�������qy���:�}ų*���@�1Xؐ%��wR)�'RY3�����\x��]�;��{&��^�J6F�H�A��P!U>�ˎǉ�T���rN{Ò6=8C�w{��odԵH�^!�9<2�$�TU��r�I?�iX>{/���r�$_cH��1-�Yo�2�!Hf���g,�Hʾ\Mz!  
KZ���{ }?��v��|�S��t�g�8k2n�Uk`rl�wp2��Y�3��t�dg�Z����+`���i������e�)]���c�V�B�x0�A�k&*�/�S��{��)S`	/��X���5��b��ߜ�S��Eli�7]�gު�평eDo+��Ѻ��L��MBJ��C�T��EY�w�Yu6�񿅗����C���x��U�p��I�Y�<�[Z���n�e�����C�Q����:���L�Y�:OS�t� �{f�(�[�Y�rm�;��S����b)��6�(��?>%Vo�0v��h4�xHPkͦ���9s_qz)U�>^����&*�%*��%%uʐ8�2Rq�x����lzQ8%�����W=������H@�¹�󌄀{v���Y�`J��:��o�N�l�O�sG����8��O��b�A�	*�2X��g0��mXlRZ}GRP5��G�w�o�^��6H׿S+Xb?dKr�����8a��;�����IB �(b��gz�!��� ,����=�p�b��a�>R%A$���iʕB�5���X,�~�#MJ���m��3��U�H}Ŷh�V���V۵=�0�N#FD�9���^
M�LG�%R�'@��6dҘ r�P��t}�o"���d>m��[�2h�-�=�M�9�ˡ�ia�bl��!��S��]d^�2m�~b\I%8�M/�}��4��J��M��Ũ@'�ݾ�o8��"�.A���IX4`D�ı��4@�Y�m�,"�u2�|�G_ڴNV9� �TP���R$p�������Gv8�"J�fm�b�����Q�{L�T1���Ģ�5��,�aܘ�o���<l�(p�������3jK��/��pk��޿����Q�S#�[mp���}<��`޺�/�5z���E�2>�ԨJJ��ÓJ\8ܜG3mQ=U������c�gFm��l��b?�����	�-���x�"\����Bz*�;���={{�J����Z]��w)�c��c-HV!������zP��9��Kŷvk"�t����Ey�sDQ������^�#��4q�n��k�$c����t��R���OP-\ �H��@&`#g?�.�EȮ2�ǽe�e��S�̼v�XȬ\(���"�=R/���at?vW7��c�3T�#&��sK8�G�VC�����=[�:ȵ]=���8�� �(R�Uˋ�'pS9l��v�Ξ���n��R���j�'�p�:�ڿ�=q���˳a��$Q��w�O�p�[s�۔��lc>nnۥ��9j؝LX6ĖѺ�{QJA�Bw��a�zȅf�R#����k�OI]Ϛ�s�$���*�uX������ڿ�&����옶fǲ�T�t1��w�C��n����RCv%�(�ee�\���g������y�H7�w�ܩ]�b��+`�o���1��ހY�C�V��.��Ӽ[@��b��:�S��������̼4��A%j!wmG/���3Ū����R{/�nHg��E�`�0���HJ"����'%9��?���T�V�� ����Zэ�۸~R������b��)���S�q<a-O�3S�G���������[ꁃb�ؗ[�@$�-�������:%��1$�x�wD�ߴ�_���U"���r�B|r���(�J"NKp�C,��msfw9(���P{���2@�ݮ�x�kQ�
��$��ӥ�6���<)DbVT��gq������z��b߈�-]C �j9o�n��E,B�F�X�}��ê,\�����rP��c���H ��%�)�u��\�]bY�f�Y]n����4����#S����C� M)������J	Agm�g#ϔ��7i~�+Z�s<:uQw��яA.`c������)4���8�E�Z�hDȄ��"���S��1!�i��>A���͔���	L? �k�-��,�=̀��|W�m�A�=<��+�pd����%VY�e�fz#�mZQ�dz�q�e�W��d�y��<G�E]�|~�\����T_�r�].(��Pj�2��4-��/�1��:>9~�L�F�(����m~W�EN6<\�5S�69�7 (���~=Ew_*���n�+�����f/�@��ጓ9|���	�z�J����j�f��_�(B�х�g����ǩ�#���ZF���x�F����C�T�B�۫�*�Z�`��!FN;Z%�>���Txi@����j����Fq2��r,_��Σ��������B[yyv�*f.����+��� v�>�tQ��:��կ5BZF*%����>ߨ�����-�{@ FYX�W���N��EvLx�@�d�Nz��i,P�p����L*��!t�b�JXl���;���E�_&H�`é�訸 Q�'V<[{��{�[qܚ�i���ݒ����>�jC����+'���e�Z��G4\kl��ʯ��t�������r<�d����ӛ��9��aHRL��bʜ}��x>W����cm@U 9}�7K謇�9�ōo��yl��ik�E��I��(�D*`��E)�,\8#4�7˪�pE{�W��X��jJ�5���o��Bb79�]L4��x�4(?/Q���0h�yB�1F��,�H'��x�����n
�l3�v�w�x��(_��y��Fv\��b*�=ş�E��Eb����*�je��\����7�q^)��[�S��[��P�91�t 68�-�m��.���um]�-��wml�Iwȋ{ ��J��4��T6�}�=�*Ώ�����O{�n���mR�&��b��|Q$N��Y"�}�X�'�
Y�S�G�j���%�:۞50{�<j~�e��;�>!�6�:M�%-�U��k[�P�v�R���4l_H�֕dMx�!ǻ(S4�"�?�K��� ͑��x����������2��\I��ۂ#-�"̜K�Q�XH���z��쨂g��βf����^��:I��3�>xS�������W�x	�=#\,�a�P�;74�7�ZDi��A-��&e+L(<���==&8
�C�ڀ�[Ѵh$7w1��ߔx�JN����5���#��r�#�>"�Iz㸄���r�"N�ӗ�b������܍q

m�%�u����4;�B�������QF�fls(�B-S�j>��ՔT��!��&�~N��̦�C|UiR�,��~�Sr�u���_��3��}��+��Ts��_A�2*N�6H�F�z�]�DV�-��:�%z��j!5sP��'�zo��	���j�e��5ɟbi�H炸�<��Gq�A_=C�$!��q\°������>�Ei�7���>�n����^�b�2���r,彩Xǻ[�_���W�QPF6��H�����*��rE
<g����]�-��Y�o��$�������ؒ�O�hO�J�����7Q������8��q�53W�S��t d<� 	�3��?�5���h��S:�\��o�S��ȖC�-��@�/E�,���C����c=�^sn������҂�*i;g��ӑ�G��=
�~ʭ�(aP:VB#V`���]���g��r���\��x��"�\�������wWV:���ٯ���8� �e���SN3����\C��[^G���^SY�a�D@˥�����ёW�%n�d�0����?eP﮵��AGY�juF4��8V�q�<-;�NJى��W�`S���=��xq�3:�$=�ssj���@b�������5*\U<:��jr�P<BW` �����	��ת&L0�\ԣp$�3�T<~�XU��)^7D;�S�[*�_���bcG"���6�>���l���lL�L�Q�Ȋu+�º��������w��U�=9!+�Hu�ƀ�|�mtJ�ϩ?��ht��c�Ԡ@������((ۜg��ɂ�QE-��o+���z�x�s͛i٦�H�>�U.�Z�tZ�>�iTO���R�.�~����$�o(��������-s�OT�s�S����_�s<�T���1%�D���q��~�3�����Ө���5��>����k#�<c�L<���lѪ���̵
1����BP��%�s�'�iC�S�^�����l�N�N��i�L����KDH� _����������Q�u͙2�=dZɿ�W�Ͼ�}���t+xR �5�b��P�9�!�D��,��L�
��j�%�L�p��f��w�<2�D�+Ғ����G�Ti@�+�g�B(���gg`�Gq>.w���Y8_]�r��{I�ڛYXQ��cpZ�[!����H�ڂԹ�2�� σ�/���ܚ�C��N�Z)+0� \<+ᠬT3�Ҥ33���D����g��*�#3Qٜ&�\ali��F�!^"%«bc��V !Fh�^{o(b�M$7���ŻI,�+�-��P�I�Zp$x�0-0�Ux�j߫�9�k��q�q��4�xp�$�o˧ ���:2���_����߂��|I�E����f�BM8�\��8�Į�7�Ӳ4�x���U�Z�<)�K�2�x��9� � Wl���3�9S��佘mZ9bB�Դ	~Y�b9�,���K�hҎ1ʘ����������NYI��a-�������1ؘay����1�D���DCEI��[U���9gZ�r]�t�!^d.x��������n�l��bw��E��3�N�y����wǃ����5�esƸ~��t������o�@�UZs��R��+b�ܑ�Bi���G�p��x4[q���yUIP����JW�����SôS��&����(t�쮊Spn��+y(|�W*�o j=�s��/�Y��/�����ܫ����t����C~�(��L�ЖF�1�#�~8U�P&�ŋ#�y+NL��V��x�ؘ_Fzզ�6�Ѿ8J<�c�+B�?,&Ξ��hv1����֔�
my4SiΧ����l�GL3 1��x�i���+h&�g��{��p��94�}��sxp;�0q��{�T&e{�+���l���j���@����d0+.��|G�MKdz��v�q������q�����p�n��*��������J�|Qq�Py2���CE�N3Ӵ&#�hk9td^�#3�`�k��6ū�#�w}4sD��� �m�|1e�l���<����}="s+fŅ�� �	HH��#���[G���>��RjPǹ�Ы �2��f�?���m��	�p�
�"�.ի�h���<5;WX,ﻜ��W�Ety��X�6�
';=��`*�Rk��@|HS�.�L��M�.�ܨa�'��Y�J��w��4%fRi��K�a��5dZ��{�^�Z>*`��W�\�pN��5�p�I��D:�3���Q�e�uWS��.���(6=^OFV�� %*<s��`���Q��]pIy���fr*��>vmӮ;�J��qA�������a�Y˵P�f�7Q��M�dtyr���h1; Y�-��J^�>[�rh�w>ђ�dy*��N��a$j.pְ��K͆'e9c�yTx����q�^Mf�S�D2�#�!>Q>�S���8�F��n	􄲏f���r�7GVu
��4��Q�9�=f���(�c��t��ix��Ym=!��w4k�Ξf����Jp�܃V�z��������v<��O�8*��r��-�=�IK�|�wx~-�kw��c��ࠧ��G�(���ό=�����+v���R�}!�c
I�׷B��"�>��(�h���8���+3�W�Pɺ2��TO^�$�~��R��J�鹎��L�7D_���]��De�B�D�����ؙ�	���$p	�
k�O��N�'Mu6��i�Ԫg�('%5*�8Wh�Qq]���j1^��.m�z��>Z7�Yg�E9�)�7
��1�A�F�,9R������o�\;N��T�*�
Z� (m���T]��*��4�ܵ����m���{K�ڨ߮͏��?�$�@p>�����!�H��;�H�
���ЈV�	i�Y� ڜRK�p��^*UC��ñ�)炼ㇷ-�-	w¶.Ow��/U��-�����Ksƞ4O�!�VV�C�7����I�c
�f&�E���$���ϓ;�&�n��%��cvc��$"�$�W�k8�h� `k1��K���uhH�9�x纡u���,�t�j�T���/����6\>�9�q��7$��N`A{�e����)�gl
���p��	ne[�&�N�
�1~nBy��_�{_i�tW��>	�hbpgS�ivY�&�9��}@�6F&�G;�|�j�{Z-�Cd��L>�ז��1o5Q>5?"�2�M�ƪn,�j�♱����������������p��է�E]1���D��
�uv#����̴�kM^��6���óU����#��8bH#�u���G�/�����G�,��z�|���#V��ti��X�-(�.�����͵`������>�)wOwf��\~E8�B����%$u6N��,j����q�ĶզNB�M��`_j8+�1/�f>dvk �F�dg0k�^s���fp,��H\Y#o�G����i��hF=��ؒ���m1�%��ּ���A|���#y���g�Bu+T���̼(��Z�x����%&�r���(Q�X���b1^��J2;z����)ds�䲂gFւR��v�y��*4n*�hM2i(�=�L�L�ǂ�zp��؆�2��=�@�uj"��9`�ɢ
�ߠm�NY�`Z� ߱�l�۱���M��9��c�D;�� Y1������1����%Uj�M��X�fd����4�qp�Ő�T�_� 7á\�о�/?���9��:����qHL}l[f�Ț}�����ܫ��u��i�F>�mje���M4��d��Y�J �a�F�d5w�����E�Utg.��2�����@�����ޤ1˻���Y�#I�o�KD���T3�{Lֶ\\�P�z
��KI������^�22ūj]Ɓ���e�+Z��E�5L[�-�Bƻ)��פ��ooY�����h�f� CK�
�P�4ahK�����K���~kʶ�r��N/񶅯Uw��C3[��f�yP6�N���Y��7�&��-��A���=�+�W�R�+�����s�?=X�!�{G����\&>1�"���T|����?�28��jF?��G^��4�p�a]�s�첑&��b\�;�gi���/���uk-��~w�g��f��2���nI�T>2#mu"v��9qx[5z7����wXD{e6;��$iyxY{�`�?�ā���!���rɳa�'�������"a�&�]����r&���j��GD)��w���U�p�W���g$���W��*-��A��J�����|Ml4R����Gi�޽���28qg}t�a>�=Ù	�vU�+V MC{�QF�ub 8~��y}�>%3C8�_VV�Va�@p�ښ������z�%6���j�s�S}g���,����`�@͛��43UB���>Ӭ�둉�c�(���*6\��p��q뵤�p�X0PBV�-�{�X���Xo��R�g�Z�J�=+@�1�I�X=� ۉ����-ɡ����vt]�S�dO`vk��^�M�V����I��v����h��5�G�/k����# �Z�fR�.��ݓ�<��u�b.�e �=Y��AU�g��a_z;��#wś��_@��lJ����m�S�>�a0�)��oHF̐L^����$����	��3Z�0.f���3�s[g[�L���6��N�~O>��e�풽�(j1,`��]`�=?�aij�+�D=Ee);"��!΁s��`��d�F�f��<�Q0@�l�P{����if��X�,O���9�I�@t����-ɷ�bU{p>�l&��ME�ε�a��Bd+�T�U�O�y�VUg�hDa"{K��0�펼4�S^�YL��1�L�w=�j�� �K�}��'9Ѐ�lgm�W������{��D\�f�C$�^�F�5����c �I�n���+��9�-���U+�����aAX���(6�a���-�LD�)B�B9 ��Ѭ��k��3<�H�����������4S����,�bzA���s��"	s����b0�����=-�1�[����6����y���X��m@�j+���W?O�)��Lʒw����΁l$H��peZ-qx^dp�T���T�>��k�����,���7��慎U$)��&כ��[k��^CmNp�'My]K��v�w��	��~'2d���^�'(r(@�#� �cP�z�h��p"c��-��7.�}+��&�<�Mi��zTcf=3�r�_ν�<vƘG��S�";��f�0�\
*��r� ��/������2��T���G��ޔt�G<3y����l}_����}��P�2Dz[���\��%�6�y2��2�ac��3v+5��o�)�'��k�ݘ�t	H�Z~��|���cжRv�:�j��&�Bz��S.񃔺7���53N_	�a�(Tgjt7ܗ�rtE�z�X�<8I���'��Kz��#\��:W��>�l����WtSwH�ʤz��`����{b*�͍�(-�z�Y��D8�����?B������x���7+y�p͕0"(�yv/�A��`���`�D���
>n�q]�0�N���r@`/hrM{|aE3㒢h�����V�q�gr){����폿���|�XBQ+�f�E�����o�3+�Y�-��CE��k��}l��B!p�ƣ.3��Mu�F�L �)]��/����Z5؂� � ����kT*
v�rU�}�����W�S�D��Y���� �g�e�!PԤ�%���(�K'����"�_cHxG��=�	 s��E�oi����2>$Y.�x�?/J@=O:�>a�'��\����wK�rG�F�&��O^̉~�kw��V� ����m�L�<�ͅD �k	9�L��ea�#����H����
n���x�:e9�죤ᰜ�B3���̭���䍸ݷr�vk�C:��w�پ�����̛])S���]J���Иg���X����b���
3q~<�ϱ�k�RYI�z _����9Yx�4��jZ}y��T&�7�᠜�f��8�=�g�|��fq�%�m������C�;͑W���5+췫����y��߭
S`�*�������)���m���7JH�b��;~`�qg��!���ю*@OX�}؏�aHu{9��]�nk
�|6��G�i��[����'�<�O�\{M?G�8=��=L��ͽ��7�tF�QN�>��&�#/i�%p��4V}��Q�!P�c�@�e`��?�=��:��Pq��ϓ�8~�[�,3��ُ������Y��K�6����}me�A,'ŕ��B�eﲼ,!�*�3΂�AY�wL�&�����^-�w�[���\_[X�0̬�L~m3)��1ۛ%��+�HfwQ62�=:���!�+�)���.��v�=��:|�������d�dO8	���澭���ѯ����b�2Y��~�bv|a>S����5S�j=cR�˷CZl�OXݴ�w�_��[���|t��;	a���{�vbm_� �~5�e���W�����t�Rj~����1�L������/��Fަ�ִ5_�@�7r<�P�q�������҅� �Y�_)��(�S$�WTAZːY��	6U�y��	8�ݹ�\d����Ubȣqhs�w+����_e+��Z1���3$�@�-�JN�\p������wW�0:����M��Mߏ�v����}�!ߥs`<��)P�8,��N�G�&� Z�n�����?*���)6~��+
wHW�BL��l(��!�K���k��,RB���3��8N9�F8�%8��{������U%j�r��`��u(��`ƥ�̱X 	/���M�_�ԴE� d-�v�{�D�`��AK6#��4�6���g&J���341��G$�fCUt��݌��.$�N�>D+���V�<L��8x�U�����}�-���I#��ovy�
�a�xn�\���� ��_�P�J��<7�G͋q���5�؆ɨ���[�te{o#ӟN�V���z�c��Յr�}�v	���q��P�D�rG�+��y^12��I������S ���!i��2��[չ�Pغ~޸*D����#o_�挰UaBfJNW�}�P���7�3$Ds2O���S�"T���%�%zX���+�2��SH/vC}s�7�06��\�t�j��3&p�23:\�u%�V$�u��PJP-\��C���]�XW����N����kʦ
� $�L�Wa/�Xn��gN
���
����$L��[S�*T��wy��%��	�/�l9ӆ����#�4g`c�e�N����G�u�>h�E-� ~�c�^��]�Vx6p��,~vpо00��(�e[r��mC\�3��Ρ��L��������wnwR��M-��7�r?&����چd��6{B�0��9�f"�
���:sy4'N��ڎ�iI�Lmcx j�L�QXϴ0U��x�@��=�ަ��^����*�9�2�
���� ���)�;���;{>� i��x���SZBM=�U�r��.�t���R��Z]�euO�ι�4�bN
 ��!�+�Fs4R�8�ɓ*yh0����Bp�FO�l���F+Ǐ���f{z� b��'�*��\�}��Cޱ�l�8�	�:��l�ZĬ�p����o��F�~����YI[I[�3��~���šSah�7�ZW+ԯz�4)�0�\мS8��Vll�f���������]��I�(OY ɇU �)���+��͌?U� �Da0H2{6R<Y���z`�e?/�)b�	3�&DcĒ�K�D�*�����E�cגO[^�GoW��I�NexL݇K�!�}�wYN\В'�F�-���H�	�f/�}e�tm���eK�a���pMo%o	�T
SZ���g�ꏍ8w�����������.Ԣ���<٥3��,\���8)j��:�Z�IpEϰOS�0� ��Ʊ��kT�ķ	IpD!t)o�>J�E�@�O��}�s��@b�v�C0�OOt��h�����k�&+��h�l����
>X]���~ZK�r�_�ӷD~���h[�
�ތ�AgT��S��f<ӊ�>�e� �q�m`���k�(8�y%~�ޡ�?����'���g��v��'0��j1������`�$$t_??��H��y@6�*5�)A��wU��~����+�p^�v�jeet�͸�{���K����f��VZ���S�W���d���n���:�ù��r	��a�z�\3r��K�Ɠ98�bo��m<$��Fm�o�����[{���7 b��p�P��Y�j+f�o-���ey�*6<O\�ꂑ��m�^`w���1�.lb,��}�p��$7��!���@���o詰Ø!����u�V��c�R�ڙ���D������Q���r	*��%�ԆM៦{�un-�<ӊ��>�k��_����׆�g���z�+f��'��;�[��� tyNB�$���a�I!_A�r��L\�L�X+�z�PF��6_�U����Z]*j�N��+�k[��.7\G�p���v��7�5ӏf�N������L?��.� K���q�\���phw��C6�߅N�>�V�NOƧ�J��d��ܢ�΄M�Y�h[�W�QOb��3,�l:pbFU�A�&+����].�,�7�7��d#చ�r�O����
���
���؟*�6��U�6�׽E���лMp6�tY+
O>�	�m����,{+�u3/|cZ��\�y�OT��0������M���
'�YC�-D�%������I�8��ANKNF��{�v�@���F�	d�cL�h``��H�8<2��L�`D
+�@����Z�	�h�lI��*�>hnl��fA��U�ýby�$Y�|�ɦM�=()�?),��`'�N�������ռ�,;��L�4U+p�>$��XѺ~!z{�s�d^�^N1�#Nm�4A��M����¬�@j�������ꦴd)���)eK�Ufؾb_���r�5$ߔZ�w�J;P���8�m�cA�(�T�U�SJ���t�#�B�c�\���H��Ao��̺�W�?4��e�ȹ�Ec��/�B�����b6m�c��d|����^�a���y���?۰��'5㿎�Z=���68��Q@��j�<� #QKr�;���&���)�k�S(�|d6?���iSTo�y�����q���2���he��tM���D��s2�@\����/��^�z	F��k��0M��9�H#jc��D��(_=D�A��p���|7�g<�k�
�iU�����NHU�⦛��M+{m��ճ&z-�r��X�(���� ^�
�$?��7�GvG���ͧ�oB���k����E�A?NW6����'�Wڣ�M����
L|>������t�����,�uU���z���$����u�J��U����x�Y��'trS�?�ͮq�*{����h��9Ԝ	�Fɕ�%`�;�4&�*��uri�qH�7�{�X=߅���p���f؀G���+���|�zp�m2Ը��`.�ԇ�s-����~�x!;]�K%�HHBn�(1dm��BEn�}�z�=�G��8��ݸ_�u��D���҈�s�.�4[��t�#��惬��+����.I��kY���Mh����GO6��-�؍�o�����T���C�4�i��0 .0��%���,p���s����ب1��,(R�P����]���/+u Ed�?��l�e�������X6��|_������	֕�3��P���+�M����� �d�+��9�Y8��V{٬��8����(=���bC�^N�(P����1륡9w٦wx���aC^pF]"�z�:h���+2�卨�#���D���u�1_�s
И�4�Z�fWF���ŕK=��!|S	:����Q2T��\��ɩ�
�GS+u?� ,l�}��3J���Q�ߙ��9�_v������b�1>J<w�æ]`t�F��UJ��}����x��z�����dk�l&�x�4��8�"e��2�/R�����>=J;!���^y�[P���@ϊ�Z')�M	ׅ��l���S�u�}��q�����A�m������������To'�n�U��2�o�Kﴖ�[��=�� ���w�a��@&�K�IF>�|�LWo�^���\EMn�c�?�Q��^���@���vgq��dS<0���ȳ`{����׽��u�@�u��rt��˟��s-:�c�pme�k�}�^9w�� GA�t�铊�N9oV�աד�Lƥ}JHw� �}ݭ�\v��3�$�k��G����������=�,��YK�������:Ű=�%���x���D���	Տ�q���O�q� F*�-ϸv<��2��k9(��D�f]���bH�"}���m�F%��*k�8�nZ�����%m���?��z�b�M�C�!�ݼ�K^ �mI�n�8��fh@�2�{Зg��>�Cb���r�ɀrR ?Y,�5�i���]�L�n|����WQ	i��S��N�'�T#j]O�܄���\  =���~]7J���^��gO�P'��zc h�Y
d�tz�~M�tn^jɠ߽��e�J5b k
G@�$�+6%�`��b���p�4�u��64F��mm상DHqaP+e5h�%<*��%@7���PJMn��^���-C&�-ԍ��l�X݅	�
���/�s�=V�OX��v���ئ�K�1Qh��S9��6HzQmx��M�0/�����7>
��WK�d	���6������O*�Ե[�%;��B����(�F�-�h;��3�����r1;HM���rt�`�#Y��4�N�˿�-�ض�>:�{�4I�Ͷn��-��L-���X5�E�%.JXG��A����U����
�p4-.\@�J��xI��0�c� 4�R�Xuz����_������H�O���d�0wu����D�h�h�졣(H�Y�o��5ִ5/
���X�(
#̞4�kx+!�����������:b�)�{�	v,�>�{�s7_(L�#�s="��9˅�uTPǧ�\����5�R���9���'��E���}��⡻�i�W�e_ �.�Οp�� ý����0����s��������. �P�?�Ƕ���q!�[�˥�x��Nn�����_��w̪�Wz�! �:��v�el� VM)4%�n��}ѭ�q�8xa���4����%�ͮ�ߐQ���dT�#i��sFM�:��M��	�����C�������c�� ���E� ��Z�ӹ|?�p����/��ʹ��"�m��� Ip�Y��{3ΫRE0fϚ�ApF� ���:� �H/�ve�w¯~��j����u/���jVC����N�tA5�GM����F�g1��V!�4��8�<e�땿'�����)�T����4�d'3��q��$��S�j���yy��|�.~i��;W�-�� LO�8���F�C�����x*��q?�Y�˗�K$X�w;[�8����.Q6"9����yԨN�<P�����Ƚ� 9��o�Qg�c��qD+��V+d1o�h�Eg���^Z �"ͪ0V����8����ǿ��Dc���liE�hLH:�Vo5���nJ�3)�j!j��z!����9'��|px�N��~3X��*U J�K��7q�_ǫ�p�e�#c����0�r��(Z����u�z@�dv` `�儏�uT8 n
.HO&K��/-�,�,�̒HŤ_���0f��ʱ����P\�����%��M���'?cG1o)�t�m�ؼ�B�:\����z]�:�j|imRI�L���Fl�����A��a��bd���cd���C�"�]�����R�T~��p���(�J�sl)6ۃ��H&����n��erDEa�����J��OǇJ|=/�,ʤ��k�cgF�Һ:����T�[��?7���l� ^$uO�Y#I��a�����rC�������vo�}X���Eրd@9��rS�޴��@��M��̽`\�J�(jg�Q�`F}Mv��N������;D_�ܨm1�o{����T,������ɀ9�
oA��(ۇ`��_z� /��:�N5HeZO�P�cM~��A�Yh�].��Iy@F��R?5s�����|S�A(��1�c�[�
�i2��n��q��j�6A6Uɯ6�bp| *��T6Bd��=��y� �f��YӕU�e6y��E�����lr5����.�R�59�U9Cl6/#�zk�bxA4^8�L�a�Yzŷ99�3p|$��d��.��D_��@��:�#��@��u?sa��E��@���3Z�vG:�c��CzLދ��mY�3��$m��.I[&u�)�_iȁ��?����*~(����,t��'t��d;���2������⣡�Gd�A�;<��4�ۓ9�Zΰ��5祪�����$��*������h�ԬB᫮t�	垛�U�r�*���s#lTh�vVb��9����:��&G)u�x~���Q#�S�ʑ#�S�'��d���?�#B`�� �l\�2�I�
7�TFƌwjܐ|�+�q��������lo���<j�"�	�ߤ|�j��dP� s^`�hؽ�dUxRm؇�������mR��׈[%��Q��
���5�O뀧����W�j��BҜ�PK���˝���ճ����>õ��&�/���0]][~9 �Ҕ�H:�� �1����^~D�#nk�
�b�`�^���#�q��1�}2�-0y���f��<x8Z5�Ut7��:`�������HW#8�"iN�`S�ێ%1-e�&'��Ҕs�2s���s6ք��2�0����ҏo�)�8��H;��e(qnII���^�[�vV�u�B�8
��P�ǃ��c]B��rb������O��ٰ�~���	�<�x}��DJ�c�P.���r�:��60.�N�i����5��w�h��W=�&�y��t> �m	ʗi�%>�>D+�j_�y@%����7���֠�?82H�$x ��\��UҦ]����?TM/A�u ��c�U�dI��@�O��5-ԑ��#���af�::��҃&�n�oI��8jQb�u��T�� 7lS�g�^�G N=���&�93���;��I,n�%��yq��֨$�p}��1�h�1,<xCѠÞ�����μ��������Db�y�*ݟv���n����CS��gx)�>"BeQe{@e	Pf	U 83ђ(n�٩�襀���g�-�rZ�F9֦�;��l��+;'x`�%h|<�D�ey��+|�֊�w��Z��l����\�H=��;D;�V��(�]<L��!�Ǳ���� , ���miibT�<�1���յ!����(1X���8~l3S@��M2N��2Q{!�9"��yLJ��U�l}�'����+��Ç���wY8�!�Ѐ�+og�qI���)���ϊ?��o�i�&|z��6�*Yk�K'i�Or�t(�2�c��d/���ט�o�A�*6����?�=� 2�F��#�$�@���˟���%���m�>v�8��d�WK�X�a�y7�G\@���pW����2��k,�c5�]�Rm�=�G����R�,kԼx{�<l_i�y�<?P��nU���0 -�c��������� F�x�h� w �&�:m��d3/7��dLpn�\O��+�bh\k{�w�⊱������A]�翖Լ���U����b��Ygq6�?��p�梫{ �o����j��C�9Ruͼɸ����Ϝ���)7���;� ���Y�7���b<�|��F��J7���A>��xy,}/N�	13U�"��;�mM+�+��%fC���Q��a�\�ԡ�qR�p��}���(VF3��: #l�efO��乭0Q�n�z�_�$0ߤ�O�U��>biX<D�;�|)'O��^�P$�t� ���Sh'�V��>��CRlb���ذ�V�������� �h{i�p���v��ځ�!�&E'ʌN�%h�uWp�A4c��w"q��%y����-/�Ԛ�٥�bIP��n#��gN �"iR�"���qo��� ����q�N�Oe��(2"-`Z��qZl1�p_"x&M�}����`BJ�d��^<��+2�^��	Yi���7����iܖ/���p	�}���m��#�ҫL	)ߣ����y1���W�����ӫ�=�Z�$�ַ�Z��ٜ�RA�̃�Q��S�[���P����?�g��Q1�"�W�}{)�D:�� T���O�-l��5��U���2x���q@�Nf�E+C�B�H�_�7����F��\}�0�V��/t*�O�����7[���ouU��y<�p����0 f��pF�G��s��i���#�Z�Ш��A�!�ĭb���~� ��(��"�W�lU���߲�}�P��M� t	�a{�ޔ�zs��	�� ��=��zΩ�V �QO��C��L@����nr�w1���?$yad��2��\^bv�ݝ(�E��ָ�Z�g��Ϟ��/Ǌ��c�{�G!�h����e�h�u�!Z��_+gj��5s�:xg>�k���� r�pp��p������9$<bT�c����L(�k	��T�?���7M�����<�o,���z��x�I$ã�>&�hN������(zη=mA\�xt���a}�uH�+��@��
J*e� U�u �F���e�Z����U#F�:����F�s�F?��58)���L}�m�i�r�w���e?.|nUF����g���5��j]�QXj�j1t[�ER�������/2�G>����(7vl��Ze���˷/�z��d.��}ޯ\uÎ�,tc|�~��.�'�l�����(ּ�[5ܜ�zo�c�-�
1/6���%&f^����%h�;��	�1�����j��s2OJ&.Św�R
/����{��%�#������"a�T�Ֆ	؂>���̯T��b�Fm�)=S]��Cf���m����9Q*;�6��>͕L�$�.+��h�:�f��)�����[�dK�K A!�h�g7}��ꁕ�c�F�A��~0X4��t����Y��IP���S��k������ȫ+���dZ��6{UW���۶.{������!;�Co��7Lv�������cT���}8��l�"��Բ=s�@~��դ-�l�dC|��Z�:,M��E{�Qg����qBش�o�2Y��.l�+ZpF^/q[ќ��g�'�Ԇ���v�4 ����w�z��zz�eh��T���*�)t��[#�ne"�a(�� ��47���p�6C����i	!�U+JiwfIVC���1F('R�֣�s3�_d�0mwr��?�ӥ@���(�M��*�X��З2g-�#�Ǽ)��g~L	:�҆��T%����>�DS� t
��cB�Q� �Z�PcV��[�Ҽq��܂Ov$f����,1��U��Յ!�Z鯜�6��~�^q���d+5��;�T6tg��EOi��j����M�NJ�*S*Du��}
��pe�(���[>�3�jJ.�|����Cj���;�>��||����<����5<b�AO���&�TfW��0���i"���:�j �;&J� ���X��>��"���rbl�.-�B v/��|��ަ�FS����Im�J�ۏ���-jP��%�_͑KôO���N�ò�>�_�O��&�kņ!{�Sŭ�X��ʵ@���<���x�������$s�[%Ք�\"����!v7Yg]>��FLM�A^���{ֿW�X�0�Av��tt�3�zl,N����
iM$�$c�}���
�4�N_�:��ge���f���%����q?�f���6����F]�t��Ѳ��ft�u�����)�<�Ͼb�R��\�������H`��\�=7j5�}*˜܊}��3��f�R�9U�g�]q��͑��4�����,֥�{0�G��LV��-�%
�yE���V��$C�^P�[�00d1�7(W��r��qY�T�0�W�(���c%T�JЌT��k�~��M{���I�-d���u����B�ݶI��C�G�Z�����p���<���y��uHغ�M��8�漀�1���E�����/P�bV�x
"Л��r� r��1����+�b(?�	���|^Ud������ylM6#^+[�ǚ����������&�}F�E!m����3ҕ|]����)e�˹"l5�e���7�$�ǎ�}�� �p�U'���{��8�˦��5T������A4�Rs. ����޶����!���{��y4��NTdUM';"��9Zj~�>lgR������y�Pu�q�o6ny���`䆞1K��jz� �Cs�I|55���}�
��(HZ��h}K}���>�������y�� �"�z�GjeA���q�I����;��3c��X�>�_�j�}.!�Gq�>7)Y D�n�Q��1p[v\Plk�F���R�����4h�$g�v��`WB�:Jb}����7�4W�2Cǧ��!�K`N����Z�rH��Y���`7n�C�OJ���^l���N�#�P�`M�=����h��lϛ�S��/��JF-��p}�Υ�?���>�3k�_Xa�uΌ��O�@��Ȟ���@�9���d����LD�Ѽ7�i�*/�L�!�Ĕ���T���Q p��yܮNZF5��@�2=N����h��xC�ϣ��eE�����2uw�ńt�b��Mcjh��9�����r+�Spn��o�l���3�������hw�K�(9�e��p�}c8���*Q��۱���r
�`��h���4�19�Jѐ��)��f�%�;��ȅ�����ɯؙ�2�'@ �P\�&A��U����j𣞛2U��J���W`*�����j�ժ��#|Z�Jp�N#����x����_TtX[�C�K9��5�=�˾�,<�Bf�+��G�QqJp��\�6����q:��\��r58���Y�7��GWJ�~	�w��(sBSY��A� �B�:���Ha�~� ;A�7��n� 
����J6YM��4c�j��):؃Ƃ`�w���.����=ԛ�U���.C\�Ͳ��m��&(]\/��>M[`�.��r$ַ�Tg0ʹA�UZ<�C�<xT09��N����ac4J����H�0⩶��L�=Gr�'z�^0vqE}N�������WsXf�%��`h�D*���~��	_<�ݰ�v�=t�i~�~�������[2z3nz&m��ǀ�+ �o�HVkaa�����@�%_׷�ib�΂
��!�;�<z�����PsA+`�=��ͽ/A0Ƥ���WKxv3�?z2 Beޠ�{�v��mv��/��ERz��~K+c�[����������À���a��z����a�P��R^w�U�����QY SY��2�F0{A��V�kp7C�Ԗk�����3C�v�Ә�6hh��ƅIQUl�rs �Le�$1�b���4